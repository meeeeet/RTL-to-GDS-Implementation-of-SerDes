interface if_serdes(input clk,en);
    
    logic [31:0] din;
    logic ld;
    logic [31:0] dout;
    logic ser_dout;

endinterface