module des (clock,
    din,
    enable,
    load,
    dout);
 input clock;
 input din;
 input enable;
 input load;
 output [31:0] dout;

 wire \DATA.din[0] ;
 wire \DATA.din[10] ;
 wire \DATA.din[11] ;
 wire \DATA.din[12] ;
 wire \DATA.din[13] ;
 wire \DATA.din[14] ;
 wire \DATA.din[15] ;
 wire \DATA.din[16] ;
 wire \DATA.din[17] ;
 wire \DATA.din[18] ;
 wire \DATA.din[19] ;
 wire \DATA.din[1] ;
 wire \DATA.din[20] ;
 wire \DATA.din[21] ;
 wire \DATA.din[22] ;
 wire \DATA.din[23] ;
 wire \DATA.din[24] ;
 wire \DATA.din[25] ;
 wire \DATA.din[26] ;
 wire \DATA.din[27] ;
 wire \DATA.din[28] ;
 wire \DATA.din[29] ;
 wire \DATA.din[2] ;
 wire \DATA.din[30] ;
 wire \DATA.din[31] ;
 wire \DATA.din[3] ;
 wire \DATA.din[4] ;
 wire \DATA.din[5] ;
 wire \DATA.din[6] ;
 wire \DATA.din[7] ;
 wire \DATA.din[8] ;
 wire \DATA.din[9] ;
 wire \DEMUX16X4.d_in ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire clknet_0_clock;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire net7;
 wire net6;
 wire _109_;
 wire net5;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire net4;
 wire _130_;
 wire net3;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire net2;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire net1;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire clknet_2_0__leaf_clock;
 wire clknet_2_1__leaf_clock;
 wire clknet_2_2__leaf_clock;
 wire clknet_2_3__leaf_clock;
 wire net73;
 wire net74;
 wire net75;

 TAPCELL_ASAP7_75t_SL PHY_8 ();
 TAPCELL_ASAP7_75t_SL PHY_7 ();
 AND2x4_ASAP7_75t_SL _173_ (.A(_032_),
    .B(_066_),
    .Y(_109_));
 TAPCELL_ASAP7_75t_SL PHY_6 ();
 INVx1_ASAP7_75t_SL _175_ (.A(net73),
    .Y(_111_));
 AND3x2_ASAP7_75t_SL _176_ (.A(net75),
    .B(_068_),
    .C(_111_),
    .Y(_112_));
 NAND2x1_ASAP7_75t_SL _177_ (.A(_109_),
    .B(_112_),
    .Y(_001_));
 INVx2_ASAP7_75t_SL _178_ (.A(_068_),
    .Y(_113_));
 AND3x2_ASAP7_75t_SL _179_ (.A(_067_),
    .B(_113_),
    .C(_033_),
    .Y(_114_));
 NAND2x1_ASAP7_75t_SL _180_ (.A(_109_),
    .B(_114_),
    .Y(_002_));
 AND3x2_ASAP7_75t_SL _181_ (.A(net75),
    .B(_113_),
    .C(_111_),
    .Y(_115_));
 NAND2x1_ASAP7_75t_SL _182_ (.A(_109_),
    .B(_115_),
    .Y(_003_));
 INVx1_ASAP7_75t_SL _183_ (.A(net75),
    .Y(_116_));
 AND3x2_ASAP7_75t_SL _184_ (.A(_116_),
    .B(net74),
    .C(net73),
    .Y(_117_));
 NAND2x1_ASAP7_75t_SL _185_ (.A(_109_),
    .B(_117_),
    .Y(_004_));
 NAND2x1_ASAP7_75t_SL _186_ (.A(_032_),
    .B(_066_),
    .Y(_118_));
 OR3x1_ASAP7_75t_SL _187_ (.A(_067_),
    .B(_113_),
    .C(_033_),
    .Y(_119_));
 OR2x2_ASAP7_75t_SL _188_ (.A(_118_),
    .B(_119_),
    .Y(_005_));
 AND3x2_ASAP7_75t_SL _189_ (.A(_116_),
    .B(_113_),
    .C(net73),
    .Y(_120_));
 NAND2x1_ASAP7_75t_SL _190_ (.A(_109_),
    .B(_120_),
    .Y(_006_));
 OR3x4_ASAP7_75t_SL _191_ (.A(_067_),
    .B(_068_),
    .C(_033_),
    .Y(_121_));
 OR2x2_ASAP7_75t_SL _192_ (.A(_118_),
    .B(_121_),
    .Y(_007_));
 INVx2_ASAP7_75t_SL _193_ (.A(_066_),
    .Y(_122_));
 AND2x4_ASAP7_75t_SL _194_ (.A(_032_),
    .B(_122_),
    .Y(_123_));
 AND3x2_ASAP7_75t_SL _195_ (.A(_067_),
    .B(_068_),
    .C(_033_),
    .Y(_124_));
 NAND2x1_ASAP7_75t_SL _196_ (.A(_123_),
    .B(_124_),
    .Y(_008_));
 NAND2x1_ASAP7_75t_SL _197_ (.A(_112_),
    .B(_123_),
    .Y(_009_));
 NAND2x1_ASAP7_75t_SL _198_ (.A(_114_),
    .B(_123_),
    .Y(_010_));
 NAND2x1_ASAP7_75t_SL _199_ (.A(_115_),
    .B(_123_),
    .Y(_011_));
 NAND2x1_ASAP7_75t_SL _200_ (.A(_117_),
    .B(_123_),
    .Y(_012_));
 INVx1_ASAP7_75t_SL _201_ (.A(_032_),
    .Y(_125_));
 OR3x1_ASAP7_75t_SL _202_ (.A(_125_),
    .B(_066_),
    .C(_119_),
    .Y(_013_));
 NAND2x1_ASAP7_75t_SL _203_ (.A(_120_),
    .B(_123_),
    .Y(_014_));
 OR3x1_ASAP7_75t_SL _204_ (.A(_125_),
    .B(_066_),
    .C(_121_),
    .Y(_015_));
 AND2x4_ASAP7_75t_SL _205_ (.A(_125_),
    .B(_066_),
    .Y(_126_));
 NAND2x1_ASAP7_75t_SL _206_ (.A(_124_),
    .B(_126_),
    .Y(_016_));
 NAND2x1_ASAP7_75t_SL _207_ (.A(_112_),
    .B(_126_),
    .Y(_017_));
 NAND2x1_ASAP7_75t_SL _208_ (.A(_114_),
    .B(_126_),
    .Y(_018_));
 NAND2x1_ASAP7_75t_SL _209_ (.A(_115_),
    .B(_126_),
    .Y(_019_));
 NAND2x1_ASAP7_75t_SL _210_ (.A(_117_),
    .B(_126_),
    .Y(_020_));
 OR3x1_ASAP7_75t_SL _211_ (.A(_032_),
    .B(_122_),
    .C(_119_),
    .Y(_021_));
 NAND2x1_ASAP7_75t_SL _212_ (.A(_120_),
    .B(_126_),
    .Y(_022_));
 OR3x1_ASAP7_75t_SL _213_ (.A(_032_),
    .B(_122_),
    .C(_121_),
    .Y(_023_));
 NOR2x2_ASAP7_75t_SL _214_ (.A(_032_),
    .B(_066_),
    .Y(_127_));
 NAND2x1_ASAP7_75t_SL _215_ (.A(_124_),
    .B(_127_),
    .Y(_024_));
 NAND2x1_ASAP7_75t_SL _216_ (.A(_112_),
    .B(_127_),
    .Y(_025_));
 NAND2x1_ASAP7_75t_SL _217_ (.A(_114_),
    .B(_127_),
    .Y(_026_));
 NAND2x1_ASAP7_75t_SL _218_ (.A(_115_),
    .B(_127_),
    .Y(_027_));
 NAND2x1_ASAP7_75t_SL _219_ (.A(_117_),
    .B(_127_),
    .Y(_028_));
 OR3x1_ASAP7_75t_SL _220_ (.A(_032_),
    .B(_066_),
    .C(_119_),
    .Y(_029_));
 NAND2x1_ASAP7_75t_SL _221_ (.A(_120_),
    .B(_127_),
    .Y(_030_));
 OR3x1_ASAP7_75t_SL _222_ (.A(_032_),
    .B(_066_),
    .C(_121_),
    .Y(_031_));
 NAND2x1_ASAP7_75t_SL _223_ (.A(_109_),
    .B(_124_),
    .Y(_000_));
 AND2x6_ASAP7_75t_SL _224_ (.A(net1),
    .B(net2),
    .Y(\DEMUX16X4.d_in ));
 BUFx4_ASAP7_75t_SL clkbuf_0_clock (.A(clock),
    .Y(clknet_0_clock));
 INVx1_ASAP7_75t_SL _226_ (.A(_034_),
    .Y(net28));
 INVx1_ASAP7_75t_SL _227_ (.A(_035_),
    .Y(net27));
 INVx1_ASAP7_75t_SL _228_ (.A(_036_),
    .Y(net25));
 INVx1_ASAP7_75t_SL _229_ (.A(_037_),
    .Y(net24));
 INVx1_ASAP7_75t_SL _230_ (.A(_038_),
    .Y(net23));
 INVx1_ASAP7_75t_SL _231_ (.A(_039_),
    .Y(net22));
 INVx1_ASAP7_75t_SL _232_ (.A(_040_),
    .Y(net21));
 INVx1_ASAP7_75t_SL _233_ (.A(_041_),
    .Y(net20));
 INVx1_ASAP7_75t_SL _234_ (.A(_042_),
    .Y(net19));
 INVx1_ASAP7_75t_SL _235_ (.A(_043_),
    .Y(net18));
 INVx1_ASAP7_75t_SL _236_ (.A(_044_),
    .Y(net17));
 INVx1_ASAP7_75t_SL _237_ (.A(_045_),
    .Y(net16));
 INVx1_ASAP7_75t_SL _238_ (.A(_046_),
    .Y(net14));
 INVx1_ASAP7_75t_SL _239_ (.A(_047_),
    .Y(net13));
 INVx1_ASAP7_75t_SL _240_ (.A(_048_),
    .Y(net12));
 INVx1_ASAP7_75t_SL _241_ (.A(_049_),
    .Y(net11));
 INVx1_ASAP7_75t_SL _242_ (.A(_050_),
    .Y(net10));
 INVx1_ASAP7_75t_SL _243_ (.A(_051_),
    .Y(net9));
 INVx1_ASAP7_75t_SL _244_ (.A(_052_),
    .Y(net8));
 INVx1_ASAP7_75t_SL _245_ (.A(_053_),
    .Y(net7));
 INVx1_ASAP7_75t_SL _246_ (.A(_054_),
    .Y(net6));
 INVx1_ASAP7_75t_SL _247_ (.A(_055_),
    .Y(net5));
 INVx1_ASAP7_75t_SL _248_ (.A(_056_),
    .Y(net35));
 INVx1_ASAP7_75t_SL _249_ (.A(_057_),
    .Y(net34));
 INVx1_ASAP7_75t_SL _250_ (.A(_058_),
    .Y(net33));
 INVx1_ASAP7_75t_SL _251_ (.A(_059_),
    .Y(net32));
 INVx1_ASAP7_75t_SL _252_ (.A(_060_),
    .Y(net31));
 INVx1_ASAP7_75t_SL _253_ (.A(_061_),
    .Y(net30));
 INVx1_ASAP7_75t_SL _254_ (.A(_062_),
    .Y(net29));
 INVx1_ASAP7_75t_SL _255_ (.A(_063_),
    .Y(net26));
 INVx1_ASAP7_75t_SL _256_ (.A(_064_),
    .Y(net15));
 INVx1_ASAP7_75t_SL _257_ (.A(_065_),
    .Y(net4));
 CKINVDCx20_ASAP7_75t_SL _258_ (.A(net3),
    .Y(_128_));
 TAPCELL_ASAP7_75t_SL PHY_5 ();
 AND2x2_ASAP7_75t_SL _260_ (.A(\DATA.din[0] ),
    .B(net3),
    .Y(_130_));
 AO21x1_ASAP7_75t_SL _261_ (.A1(net4),
    .A2(_128_),
    .B(_130_),
    .Y(_075_));
 TAPCELL_ASAP7_75t_SL PHY_4 ();
 AND2x2_ASAP7_75t_SL _263_ (.A(net3),
    .B(\DATA.din[1] ),
    .Y(_132_));
 AO21x1_ASAP7_75t_SL _264_ (.A1(net15),
    .A2(_128_),
    .B(_132_),
    .Y(_076_));
 AND2x2_ASAP7_75t_SL _265_ (.A(net3),
    .B(\DATA.din[2] ),
    .Y(_133_));
 AO21x1_ASAP7_75t_SL _266_ (.A1(net26),
    .A2(_128_),
    .B(_133_),
    .Y(_077_));
 AND2x2_ASAP7_75t_SL _267_ (.A(net3),
    .B(\DATA.din[3] ),
    .Y(_134_));
 AO21x1_ASAP7_75t_SL _268_ (.A1(net29),
    .A2(_128_),
    .B(_134_),
    .Y(_078_));
 AND2x2_ASAP7_75t_SL _269_ (.A(net3),
    .B(\DATA.din[4] ),
    .Y(_135_));
 AO21x1_ASAP7_75t_SL _270_ (.A1(net30),
    .A2(_128_),
    .B(_135_),
    .Y(_079_));
 AND2x2_ASAP7_75t_SL _271_ (.A(net3),
    .B(\DATA.din[5] ),
    .Y(_136_));
 AO21x1_ASAP7_75t_SL _272_ (.A1(net31),
    .A2(_128_),
    .B(_136_),
    .Y(_080_));
 AND2x2_ASAP7_75t_SL _273_ (.A(net3),
    .B(\DATA.din[6] ),
    .Y(_137_));
 AO21x1_ASAP7_75t_SL _274_ (.A1(net32),
    .A2(_128_),
    .B(_137_),
    .Y(_081_));
 TAPCELL_ASAP7_75t_SL PHY_3 ();
 AND2x2_ASAP7_75t_SL _276_ (.A(net3),
    .B(\DATA.din[7] ),
    .Y(_139_));
 AO21x1_ASAP7_75t_SL _277_ (.A1(net33),
    .A2(_128_),
    .B(_139_),
    .Y(_082_));
 AND2x2_ASAP7_75t_SL _278_ (.A(net3),
    .B(\DATA.din[8] ),
    .Y(_140_));
 AO21x1_ASAP7_75t_SL _279_ (.A1(net34),
    .A2(_128_),
    .B(_140_),
    .Y(_083_));
 AND2x2_ASAP7_75t_SL _280_ (.A(net3),
    .B(\DATA.din[9] ),
    .Y(_141_));
 AO21x1_ASAP7_75t_SL _281_ (.A1(net35),
    .A2(_128_),
    .B(_141_),
    .Y(_084_));
 AND2x2_ASAP7_75t_SL _282_ (.A(net3),
    .B(\DATA.din[10] ),
    .Y(_142_));
 AO21x1_ASAP7_75t_SL _283_ (.A1(net5),
    .A2(_128_),
    .B(_142_),
    .Y(_085_));
 TAPCELL_ASAP7_75t_SL PHY_2 ();
 AND2x2_ASAP7_75t_SL _285_ (.A(net3),
    .B(\DATA.din[11] ),
    .Y(_144_));
 AO21x1_ASAP7_75t_SL _286_ (.A1(net6),
    .A2(_128_),
    .B(_144_),
    .Y(_086_));
 AND2x2_ASAP7_75t_SL _287_ (.A(net3),
    .B(\DATA.din[12] ),
    .Y(_145_));
 AO21x1_ASAP7_75t_SL _288_ (.A1(net7),
    .A2(_128_),
    .B(_145_),
    .Y(_087_));
 AND2x2_ASAP7_75t_SL _289_ (.A(net3),
    .B(\DATA.din[13] ),
    .Y(_146_));
 AO21x1_ASAP7_75t_SL _290_ (.A1(net8),
    .A2(_128_),
    .B(_146_),
    .Y(_088_));
 AND2x2_ASAP7_75t_SL _291_ (.A(net3),
    .B(\DATA.din[14] ),
    .Y(_147_));
 AO21x1_ASAP7_75t_SL _292_ (.A1(net9),
    .A2(_128_),
    .B(_147_),
    .Y(_089_));
 AND2x2_ASAP7_75t_SL _293_ (.A(net3),
    .B(\DATA.din[15] ),
    .Y(_148_));
 AO21x1_ASAP7_75t_SL _294_ (.A1(net10),
    .A2(_128_),
    .B(_148_),
    .Y(_090_));
 AND2x2_ASAP7_75t_SL _295_ (.A(net3),
    .B(\DATA.din[16] ),
    .Y(_149_));
 AO21x1_ASAP7_75t_SL _296_ (.A1(net11),
    .A2(_128_),
    .B(_149_),
    .Y(_091_));
 TAPCELL_ASAP7_75t_SL PHY_1 ();
 AND2x2_ASAP7_75t_SL _298_ (.A(net3),
    .B(\DATA.din[17] ),
    .Y(_151_));
 AO21x1_ASAP7_75t_SL _299_ (.A1(net12),
    .A2(_128_),
    .B(_151_),
    .Y(_092_));
 AND2x2_ASAP7_75t_SL _300_ (.A(net3),
    .B(\DATA.din[18] ),
    .Y(_152_));
 AO21x1_ASAP7_75t_SL _301_ (.A1(net13),
    .A2(_128_),
    .B(_152_),
    .Y(_093_));
 AND2x2_ASAP7_75t_SL _302_ (.A(net3),
    .B(\DATA.din[19] ),
    .Y(_153_));
 AO21x1_ASAP7_75t_SL _303_ (.A1(net14),
    .A2(_128_),
    .B(_153_),
    .Y(_094_));
 AND2x2_ASAP7_75t_SL _304_ (.A(net3),
    .B(\DATA.din[20] ),
    .Y(_154_));
 AO21x1_ASAP7_75t_SL _305_ (.A1(net16),
    .A2(_128_),
    .B(_154_),
    .Y(_095_));
 TAPCELL_ASAP7_75t_SL PHY_0 ();
 AND2x2_ASAP7_75t_SL _307_ (.A(net3),
    .B(\DATA.din[21] ),
    .Y(_156_));
 AO21x1_ASAP7_75t_SL _308_ (.A1(net17),
    .A2(_128_),
    .B(_156_),
    .Y(_096_));
 AND2x2_ASAP7_75t_SL _309_ (.A(net3),
    .B(\DATA.din[22] ),
    .Y(_157_));
 AO21x1_ASAP7_75t_SL _310_ (.A1(net18),
    .A2(_128_),
    .B(_157_),
    .Y(_097_));
 AND2x2_ASAP7_75t_SL _311_ (.A(net3),
    .B(\DATA.din[23] ),
    .Y(_158_));
 AO21x1_ASAP7_75t_SL _312_ (.A1(net19),
    .A2(_128_),
    .B(_158_),
    .Y(_098_));
 AND2x2_ASAP7_75t_SL _313_ (.A(net3),
    .B(\DATA.din[24] ),
    .Y(_159_));
 AO21x1_ASAP7_75t_SL _314_ (.A1(net20),
    .A2(_128_),
    .B(_159_),
    .Y(_099_));
 AND2x2_ASAP7_75t_SL _315_ (.A(net3),
    .B(\DATA.din[25] ),
    .Y(_160_));
 AO21x1_ASAP7_75t_SL _316_ (.A1(net21),
    .A2(_128_),
    .B(_160_),
    .Y(_100_));
 AND2x2_ASAP7_75t_SL _317_ (.A(net3),
    .B(\DATA.din[26] ),
    .Y(_161_));
 AO21x1_ASAP7_75t_SL _318_ (.A1(net22),
    .A2(_128_),
    .B(_161_),
    .Y(_101_));
 AND2x2_ASAP7_75t_SL _319_ (.A(net3),
    .B(\DATA.din[27] ),
    .Y(_162_));
 AO21x1_ASAP7_75t_SL _320_ (.A1(net23),
    .A2(_128_),
    .B(_162_),
    .Y(_102_));
 AND2x2_ASAP7_75t_SL _321_ (.A(net3),
    .B(\DATA.din[28] ),
    .Y(_163_));
 AO21x1_ASAP7_75t_SL _322_ (.A1(net24),
    .A2(_128_),
    .B(_163_),
    .Y(_103_));
 AND2x2_ASAP7_75t_SL _323_ (.A(net3),
    .B(\DATA.din[29] ),
    .Y(_164_));
 AO21x1_ASAP7_75t_SL _324_ (.A1(net25),
    .A2(_128_),
    .B(_164_),
    .Y(_104_));
 AND2x2_ASAP7_75t_SL _325_ (.A(net3),
    .B(\DATA.din[30] ),
    .Y(_165_));
 AO21x1_ASAP7_75t_SL _326_ (.A1(net27),
    .A2(_128_),
    .B(_165_),
    .Y(_105_));
 AND2x2_ASAP7_75t_SL _327_ (.A(net3),
    .B(\DATA.din[31] ),
    .Y(_166_));
 AO21x1_ASAP7_75t_SL _328_ (.A1(net28),
    .A2(_128_),
    .B(_166_),
    .Y(_106_));
 AND2x2_ASAP7_75t_SL _329_ (.A(net73),
    .B(_128_),
    .Y(_070_));
 XOR2x1_ASAP7_75t_SL _330_ (.A(net74),
    .Y(_167_),
    .B(net73));
 AND2x2_ASAP7_75t_SL _331_ (.A(_128_),
    .B(_167_),
    .Y(_071_));
 AO21x1_ASAP7_75t_SL _332_ (.A1(_113_),
    .A2(_111_),
    .B(_116_),
    .Y(_168_));
 AND3x1_ASAP7_75t_SL _333_ (.A(_128_),
    .B(_121_),
    .C(_168_),
    .Y(_072_));
 XNOR2x1_ASAP7_75t_SL _334_ (.B(_121_),
    .Y(_169_),
    .A(_122_));
 AND2x2_ASAP7_75t_SL _335_ (.A(_128_),
    .B(_169_),
    .Y(_073_));
 OAI21x1_ASAP7_75t_SL _336_ (.A1(_066_),
    .A2(_121_),
    .B(_032_),
    .Y(_170_));
 AND3x1_ASAP7_75t_SL _337_ (.A(_128_),
    .B(_031_),
    .C(_170_),
    .Y(_074_));
 DLLx1_ASAP7_75t_SL _338_ (.CLK(_013_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[13] ));
 DLLx1_ASAP7_75t_SL _339_ (.CLK(_004_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[4] ));
 DLLx1_ASAP7_75t_SL _340_ (.CLK(_010_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[10] ));
 DLLx1_ASAP7_75t_SL _341_ (.CLK(_023_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[23] ));
 DLLx1_ASAP7_75t_SL _342_ (.CLK(_003_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[3] ));
 DLLx1_ASAP7_75t_SL _343_ (.CLK(_014_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[14] ));
 DLLx1_ASAP7_75t_SL _344_ (.CLK(_019_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[19] ));
 DLLx1_ASAP7_75t_SL _345_ (.CLK(_002_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[2] ));
 DLLx1_ASAP7_75t_SL _346_ (.CLK(_024_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[24] ));
 DLLx1_ASAP7_75t_SL _347_ (.CLK(_009_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[9] ));
 DLLx1_ASAP7_75t_SL _348_ (.CLK(_001_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[1] ));
 DLLx1_ASAP7_75t_SL _349_ (.CLK(_017_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[17] ));
 DLLx1_ASAP7_75t_SL _350_ (.CLK(_025_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[25] ));
 DLLx1_ASAP7_75t_SL _351_ (.CLK(_000_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[0] ));
 DLLx1_ASAP7_75t_SL _352_ (.CLK(_012_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[12] ));
 DLLx1_ASAP7_75t_SL _353_ (.CLK(_008_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[8] ));
 DLLx1_ASAP7_75t_SL _354_ (.CLK(_026_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[26] ));
 DLLx1_ASAP7_75t_SL _355_ (.CLK(_020_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[20] ));
 DLLx1_ASAP7_75t_SL _356_ (.CLK(_016_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[16] ));
 DLLx1_ASAP7_75t_SL _357_ (.CLK(_027_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[27] ));
 DLLx1_ASAP7_75t_SL _358_ (.CLK(_007_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[7] ));
 DLLx1_ASAP7_75t_SL _359_ (.CLK(_015_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[15] ));
 DLLx1_ASAP7_75t_SL _360_ (.CLK(_028_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[28] ));
 DLLx1_ASAP7_75t_SL _361_ (.CLK(_021_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[21] ));
 DLLx1_ASAP7_75t_SL _362_ (.CLK(_006_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[6] ));
 DLLx1_ASAP7_75t_SL _363_ (.CLK(_029_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[29] ));
 DLLx1_ASAP7_75t_SL _364_ (.CLK(_011_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[11] ));
 DLLx1_ASAP7_75t_SL _365_ (.CLK(_018_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[18] ));
 DLLx1_ASAP7_75t_SL _366_ (.CLK(_030_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[30] ));
 DLLx1_ASAP7_75t_SL _367_ (.CLK(_005_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[5] ));
 DLLx1_ASAP7_75t_SL _368_ (.CLK(_022_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[22] ));
 DLLx1_ASAP7_75t_SL _369_ (.CLK(_031_),
    .D(\DEMUX16X4.d_in ),
    .Q(\DATA.din[31] ));
 DFFLQNx1_ASAP7_75t_SL _370_ (.CLK(net72),
    .D(_070_),
    .QN(_033_));
 DFFLQNx1_ASAP7_75t_SL _371_ (.CLK(net71),
    .D(_071_),
    .QN(_068_));
 DFFLQNx1_ASAP7_75t_SL _372_ (.CLK(net70),
    .D(_072_),
    .QN(_067_));
 DFFLQNx1_ASAP7_75t_SL _373_ (.CLK(net69),
    .D(_073_),
    .QN(_066_));
 DFFLQNx1_ASAP7_75t_SL _374_ (.CLK(net68),
    .D(_074_),
    .QN(_032_));
 DFFLQNx2_ASAP7_75t_SL _375_ (.QN(_065_),
    .CLK(net67),
    .D(_075_));
 DFFLQNx2_ASAP7_75t_SL _376_ (.QN(_064_),
    .CLK(net66),
    .D(_076_));
 DFFLQNx2_ASAP7_75t_SL _377_ (.QN(_063_),
    .CLK(net65),
    .D(_077_));
 DFFLQNx2_ASAP7_75t_SL _378_ (.QN(_062_),
    .CLK(net64),
    .D(_078_));
 DFFLQNx2_ASAP7_75t_SL _379_ (.QN(_061_),
    .CLK(net63),
    .D(_079_));
 DFFLQNx2_ASAP7_75t_SL _380_ (.QN(_060_),
    .CLK(net62),
    .D(_080_));
 DFFLQNx2_ASAP7_75t_SL _381_ (.QN(_059_),
    .CLK(net61),
    .D(_081_));
 DFFLQNx2_ASAP7_75t_SL _382_ (.QN(_058_),
    .CLK(net60),
    .D(_082_));
 DFFLQNx2_ASAP7_75t_SL _383_ (.QN(_057_),
    .CLK(net59),
    .D(_083_));
 DFFLQNx2_ASAP7_75t_SL _384_ (.QN(_056_),
    .CLK(net58),
    .D(_084_));
 DFFLQNx2_ASAP7_75t_SL _385_ (.QN(_055_),
    .CLK(net57),
    .D(_085_));
 DFFLQNx2_ASAP7_75t_SL _386_ (.QN(_054_),
    .CLK(net56),
    .D(_086_));
 DFFLQNx2_ASAP7_75t_SL _387_ (.QN(_053_),
    .CLK(net55),
    .D(_087_));
 DFFLQNx2_ASAP7_75t_SL _388_ (.QN(_052_),
    .CLK(net54),
    .D(_088_));
 DFFLQNx2_ASAP7_75t_SL _389_ (.QN(_051_),
    .CLK(net53),
    .D(_089_));
 DFFLQNx2_ASAP7_75t_SL _390_ (.QN(_050_),
    .CLK(net52),
    .D(_090_));
 DFFLQNx2_ASAP7_75t_SL _391_ (.QN(_049_),
    .CLK(net51),
    .D(_091_));
 DFFLQNx2_ASAP7_75t_SL _392_ (.QN(_048_),
    .CLK(net50),
    .D(_092_));
 DFFLQNx2_ASAP7_75t_SL _393_ (.QN(_047_),
    .CLK(net49),
    .D(_093_));
 DFFLQNx2_ASAP7_75t_SL _394_ (.QN(_046_),
    .CLK(net48),
    .D(_094_));
 DFFLQNx2_ASAP7_75t_SL _395_ (.QN(_045_),
    .CLK(net47),
    .D(_095_));
 DFFLQNx2_ASAP7_75t_SL _396_ (.QN(_044_),
    .CLK(net46),
    .D(_096_));
 DFFLQNx2_ASAP7_75t_SL _397_ (.QN(_043_),
    .CLK(net45),
    .D(_097_));
 DFFLQNx2_ASAP7_75t_SL _398_ (.QN(_042_),
    .CLK(net44),
    .D(_098_));
 DFFLQNx2_ASAP7_75t_SL _399_ (.QN(_041_),
    .CLK(net43),
    .D(_099_));
 DFFLQNx2_ASAP7_75t_SL _400_ (.QN(_040_),
    .CLK(net42),
    .D(_100_));
 DFFLQNx2_ASAP7_75t_SL _401_ (.QN(_039_),
    .CLK(net41),
    .D(_101_));
 DFFLQNx2_ASAP7_75t_SL _402_ (.QN(_038_),
    .CLK(net40),
    .D(_102_));
 DFFLQNx2_ASAP7_75t_SL _403_ (.QN(_037_),
    .CLK(net39),
    .D(_103_));
 DFFLQNx2_ASAP7_75t_SL _404_ (.QN(_036_),
    .CLK(net38),
    .D(_104_));
 DFFLQNx2_ASAP7_75t_SL _405_ (.QN(_035_),
    .CLK(net37),
    .D(_105_));
 DFFLQNx2_ASAP7_75t_SL _406_ (.QN(_034_),
    .CLK(net36),
    .D(_106_));
 TAPCELL_ASAP7_75t_SL PHY_9 ();
 TAPCELL_ASAP7_75t_SL PHY_10 ();
 TAPCELL_ASAP7_75t_SL PHY_11 ();
 TAPCELL_ASAP7_75t_SL PHY_12 ();
 TAPCELL_ASAP7_75t_SL PHY_13 ();
 TAPCELL_ASAP7_75t_SL PHY_14 ();
 TAPCELL_ASAP7_75t_SL PHY_15 ();
 TAPCELL_ASAP7_75t_SL PHY_16 ();
 TAPCELL_ASAP7_75t_SL PHY_17 ();
 TAPCELL_ASAP7_75t_SL PHY_18 ();
 TAPCELL_ASAP7_75t_SL PHY_19 ();
 TAPCELL_ASAP7_75t_SL PHY_20 ();
 TAPCELL_ASAP7_75t_SL PHY_21 ();
 TAPCELL_ASAP7_75t_SL PHY_22 ();
 TAPCELL_ASAP7_75t_SL PHY_23 ();
 TAPCELL_ASAP7_75t_SL PHY_24 ();
 TAPCELL_ASAP7_75t_SL PHY_25 ();
 TAPCELL_ASAP7_75t_SL PHY_26 ();
 TAPCELL_ASAP7_75t_SL PHY_27 ();
 TAPCELL_ASAP7_75t_SL PHY_28 ();
 TAPCELL_ASAP7_75t_SL PHY_29 ();
 TAPCELL_ASAP7_75t_SL PHY_30 ();
 TAPCELL_ASAP7_75t_SL PHY_31 ();
 TAPCELL_ASAP7_75t_SL PHY_32 ();
 TAPCELL_ASAP7_75t_SL PHY_33 ();
 TAPCELL_ASAP7_75t_SL PHY_34 ();
 TAPCELL_ASAP7_75t_SL PHY_35 ();
 TAPCELL_ASAP7_75t_SL PHY_36 ();
 TAPCELL_ASAP7_75t_SL PHY_37 ();
 TAPCELL_ASAP7_75t_SL PHY_38 ();
 TAPCELL_ASAP7_75t_SL PHY_39 ();
 TAPCELL_ASAP7_75t_SL PHY_40 ();
 TAPCELL_ASAP7_75t_SL PHY_41 ();
 TAPCELL_ASAP7_75t_SL PHY_42 ();
 TAPCELL_ASAP7_75t_SL PHY_43 ();
 TAPCELL_ASAP7_75t_SL PHY_44 ();
 TAPCELL_ASAP7_75t_SL PHY_45 ();
 TAPCELL_ASAP7_75t_SL PHY_46 ();
 TAPCELL_ASAP7_75t_SL PHY_47 ();
 TAPCELL_ASAP7_75t_SL PHY_48 ();
 TAPCELL_ASAP7_75t_SL PHY_49 ();
 TAPCELL_ASAP7_75t_SL PHY_50 ();
 TAPCELL_ASAP7_75t_SL PHY_51 ();
 TAPCELL_ASAP7_75t_SL PHY_52 ();
 TAPCELL_ASAP7_75t_SL PHY_53 ();
 TAPCELL_ASAP7_75t_SL PHY_54 ();
 TAPCELL_ASAP7_75t_SL PHY_55 ();
 TAPCELL_ASAP7_75t_SL PHY_56 ();
 TAPCELL_ASAP7_75t_SL PHY_57 ();
 TAPCELL_ASAP7_75t_SL PHY_58 ();
 TAPCELL_ASAP7_75t_SL PHY_59 ();
 TAPCELL_ASAP7_75t_SL PHY_60 ();
 TAPCELL_ASAP7_75t_SL PHY_61 ();
 TAPCELL_ASAP7_75t_SL PHY_62 ();
 TAPCELL_ASAP7_75t_SL PHY_63 ();
 TAPCELL_ASAP7_75t_SL PHY_64 ();
 TAPCELL_ASAP7_75t_SL PHY_65 ();
 TAPCELL_ASAP7_75t_SL PHY_66 ();
 TAPCELL_ASAP7_75t_SL PHY_67 ();
 TAPCELL_ASAP7_75t_SL PHY_68 ();
 TAPCELL_ASAP7_75t_SL PHY_69 ();
 TAPCELL_ASAP7_75t_SL PHY_70 ();
 TAPCELL_ASAP7_75t_SL PHY_71 ();
 TAPCELL_ASAP7_75t_SL PHY_72 ();
 TAPCELL_ASAP7_75t_SL PHY_73 ();
 TAPCELL_ASAP7_75t_SL PHY_74 ();
 TAPCELL_ASAP7_75t_SL PHY_75 ();
 TAPCELL_ASAP7_75t_SL PHY_76 ();
 TAPCELL_ASAP7_75t_SL PHY_77 ();
 TAPCELL_ASAP7_75t_SL PHY_78 ();
 TAPCELL_ASAP7_75t_SL PHY_79 ();
 TAPCELL_ASAP7_75t_SL PHY_80 ();
 TAPCELL_ASAP7_75t_SL PHY_81 ();
 TAPCELL_ASAP7_75t_SL PHY_82 ();
 TAPCELL_ASAP7_75t_SL PHY_83 ();
 TAPCELL_ASAP7_75t_SL PHY_84 ();
 TAPCELL_ASAP7_75t_SL PHY_85 ();
 TAPCELL_ASAP7_75t_SL PHY_86 ();
 TAPCELL_ASAP7_75t_SL PHY_87 ();
 TAPCELL_ASAP7_75t_SL PHY_88 ();
 TAPCELL_ASAP7_75t_SL PHY_89 ();
 TAPCELL_ASAP7_75t_SL PHY_90 ();
 TAPCELL_ASAP7_75t_SL PHY_91 ();
 TAPCELL_ASAP7_75t_SL PHY_92 ();
 TAPCELL_ASAP7_75t_SL PHY_93 ();
 TAPCELL_ASAP7_75t_SL PHY_94 ();
 TAPCELL_ASAP7_75t_SL PHY_95 ();
 TAPCELL_ASAP7_75t_SL PHY_96 ();
 TAPCELL_ASAP7_75t_SL PHY_97 ();
 TAPCELL_ASAP7_75t_SL PHY_98 ();
 TAPCELL_ASAP7_75t_SL PHY_99 ();
 TAPCELL_ASAP7_75t_SL PHY_100 ();
 TAPCELL_ASAP7_75t_SL PHY_101 ();
 TAPCELL_ASAP7_75t_SL PHY_102 ();
 TAPCELL_ASAP7_75t_SL PHY_103 ();
 TAPCELL_ASAP7_75t_SL PHY_104 ();
 TAPCELL_ASAP7_75t_SL PHY_105 ();
 TAPCELL_ASAP7_75t_SL PHY_106 ();
 TAPCELL_ASAP7_75t_SL PHY_107 ();
 TAPCELL_ASAP7_75t_SL PHY_108 ();
 TAPCELL_ASAP7_75t_SL PHY_109 ();
 TAPCELL_ASAP7_75t_SL PHY_110 ();
 TAPCELL_ASAP7_75t_SL PHY_111 ();
 TAPCELL_ASAP7_75t_SL PHY_112 ();
 TAPCELL_ASAP7_75t_SL PHY_113 ();
 TAPCELL_ASAP7_75t_SL PHY_114 ();
 TAPCELL_ASAP7_75t_SL PHY_115 ();
 TAPCELL_ASAP7_75t_SL PHY_116 ();
 TAPCELL_ASAP7_75t_SL PHY_117 ();
 TAPCELL_ASAP7_75t_SL PHY_118 ();
 TAPCELL_ASAP7_75t_SL PHY_119 ();
 TAPCELL_ASAP7_75t_SL PHY_120 ();
 TAPCELL_ASAP7_75t_SL PHY_121 ();
 TAPCELL_ASAP7_75t_SL PHY_122 ();
 TAPCELL_ASAP7_75t_SL PHY_123 ();
 TAPCELL_ASAP7_75t_SL PHY_124 ();
 TAPCELL_ASAP7_75t_SL PHY_125 ();
 TAPCELL_ASAP7_75t_SL PHY_126 ();
 TAPCELL_ASAP7_75t_SL PHY_127 ();
 BUFx2_ASAP7_75t_SL input1 (.A(din),
    .Y(net1));
 BUFx2_ASAP7_75t_SL input2 (.A(enable),
    .Y(net2));
 BUFx16f_ASAP7_75t_SL input3 (.A(load),
    .Y(net3));
 BUFx2_ASAP7_75t_SL output4 (.A(net4),
    .Y(dout[0]));
 BUFx2_ASAP7_75t_SL output5 (.A(net5),
    .Y(dout[10]));
 BUFx2_ASAP7_75t_SL output6 (.A(net6),
    .Y(dout[11]));
 BUFx2_ASAP7_75t_SL output7 (.A(net7),
    .Y(dout[12]));
 BUFx2_ASAP7_75t_SL output8 (.A(net8),
    .Y(dout[13]));
 BUFx2_ASAP7_75t_SL output9 (.A(net9),
    .Y(dout[14]));
 BUFx2_ASAP7_75t_SL output10 (.A(net10),
    .Y(dout[15]));
 BUFx2_ASAP7_75t_SL output11 (.A(net11),
    .Y(dout[16]));
 BUFx2_ASAP7_75t_SL output12 (.A(net12),
    .Y(dout[17]));
 BUFx2_ASAP7_75t_SL output13 (.A(net13),
    .Y(dout[18]));
 BUFx2_ASAP7_75t_SL output14 (.A(net14),
    .Y(dout[19]));
 BUFx2_ASAP7_75t_SL output15 (.A(net15),
    .Y(dout[1]));
 BUFx2_ASAP7_75t_SL output16 (.A(net16),
    .Y(dout[20]));
 BUFx2_ASAP7_75t_SL output17 (.A(net17),
    .Y(dout[21]));
 BUFx2_ASAP7_75t_SL output18 (.A(net18),
    .Y(dout[22]));
 BUFx2_ASAP7_75t_SL output19 (.A(net19),
    .Y(dout[23]));
 BUFx2_ASAP7_75t_SL output20 (.A(net20),
    .Y(dout[24]));
 BUFx2_ASAP7_75t_SL output21 (.A(net21),
    .Y(dout[25]));
 BUFx2_ASAP7_75t_SL output22 (.A(net22),
    .Y(dout[26]));
 BUFx2_ASAP7_75t_SL output23 (.A(net23),
    .Y(dout[27]));
 BUFx2_ASAP7_75t_SL output24 (.A(net24),
    .Y(dout[28]));
 BUFx2_ASAP7_75t_SL output25 (.A(net25),
    .Y(dout[29]));
 BUFx2_ASAP7_75t_SL output26 (.A(net26),
    .Y(dout[2]));
 BUFx2_ASAP7_75t_SL output27 (.A(net27),
    .Y(dout[30]));
 BUFx2_ASAP7_75t_SL output28 (.A(net28),
    .Y(dout[31]));
 BUFx2_ASAP7_75t_SL output29 (.A(net29),
    .Y(dout[3]));
 BUFx2_ASAP7_75t_SL output30 (.A(net30),
    .Y(dout[4]));
 BUFx2_ASAP7_75t_SL output31 (.A(net31),
    .Y(dout[5]));
 BUFx2_ASAP7_75t_SL output32 (.A(net32),
    .Y(dout[6]));
 BUFx2_ASAP7_75t_SL output33 (.A(net33),
    .Y(dout[7]));
 BUFx2_ASAP7_75t_SL output34 (.A(net34),
    .Y(dout[8]));
 BUFx2_ASAP7_75t_SL output35 (.A(net35),
    .Y(dout[9]));
 INVx1_ASAP7_75t_SL _225__1 (.A(clknet_2_2__leaf_clock),
    .Y(net36));
 INVx1_ASAP7_75t_SL _225__2 (.A(clknet_2_0__leaf_clock),
    .Y(net37));
 INVx1_ASAP7_75t_SL _225__3 (.A(clknet_2_2__leaf_clock),
    .Y(net38));
 INVx1_ASAP7_75t_SL _225__4 (.A(clknet_2_0__leaf_clock),
    .Y(net39));
 INVx1_ASAP7_75t_SL _225__5 (.A(clknet_2_1__leaf_clock),
    .Y(net40));
 INVx1_ASAP7_75t_SL _225__6 (.A(clknet_2_1__leaf_clock),
    .Y(net41));
 INVx1_ASAP7_75t_SL _225__7 (.A(clknet_2_1__leaf_clock),
    .Y(net42));
 INVx1_ASAP7_75t_SL _225__8 (.A(clknet_2_3__leaf_clock),
    .Y(net43));
 INVx1_ASAP7_75t_SL _225__9 (.A(clknet_2_2__leaf_clock),
    .Y(net44));
 INVx1_ASAP7_75t_SL _225__10 (.A(clknet_2_0__leaf_clock),
    .Y(net45));
 INVx1_ASAP7_75t_SL _225__11 (.A(clknet_2_3__leaf_clock),
    .Y(net46));
 INVx1_ASAP7_75t_SL _225__12 (.A(clknet_2_1__leaf_clock),
    .Y(net47));
 INVx1_ASAP7_75t_SL _225__13 (.A(clknet_2_1__leaf_clock),
    .Y(net48));
 INVx1_ASAP7_75t_SL _225__14 (.A(clknet_2_1__leaf_clock),
    .Y(net49));
 INVx1_ASAP7_75t_SL _225__15 (.A(clknet_2_3__leaf_clock),
    .Y(net50));
 INVx1_ASAP7_75t_SL _225__16 (.A(clknet_2_3__leaf_clock),
    .Y(net51));
 INVx1_ASAP7_75t_SL _225__17 (.A(clknet_2_2__leaf_clock),
    .Y(net52));
 INVx1_ASAP7_75t_SL _225__18 (.A(clknet_2_0__leaf_clock),
    .Y(net53));
 INVx1_ASAP7_75t_SL _225__19 (.A(clknet_2_3__leaf_clock),
    .Y(net54));
 INVx1_ASAP7_75t_SL _225__20 (.A(clknet_2_1__leaf_clock),
    .Y(net55));
 INVx1_ASAP7_75t_SL _225__21 (.A(clknet_2_1__leaf_clock),
    .Y(net56));
 INVx1_ASAP7_75t_SL _225__22 (.A(clknet_2_0__leaf_clock),
    .Y(net57));
 INVx1_ASAP7_75t_SL _225__23 (.A(clknet_2_3__leaf_clock),
    .Y(net58));
 INVx1_ASAP7_75t_SL _225__24 (.A(clknet_2_3__leaf_clock),
    .Y(net59));
 INVx1_ASAP7_75t_SL _225__25 (.A(clknet_2_2__leaf_clock),
    .Y(net60));
 INVx1_ASAP7_75t_SL _225__26 (.A(clknet_2_0__leaf_clock),
    .Y(net61));
 INVx1_ASAP7_75t_SL _225__27 (.A(clknet_2_2__leaf_clock),
    .Y(net62));
 INVx1_ASAP7_75t_SL _225__28 (.A(clknet_2_0__leaf_clock),
    .Y(net63));
 INVx1_ASAP7_75t_SL _225__29 (.A(clknet_2_0__leaf_clock),
    .Y(net64));
 INVx1_ASAP7_75t_SL _225__30 (.A(clknet_2_0__leaf_clock),
    .Y(net65));
 INVx1_ASAP7_75t_SL _225__31 (.A(clknet_2_2__leaf_clock),
    .Y(net66));
 INVx1_ASAP7_75t_SL _225__32 (.A(clknet_2_2__leaf_clock),
    .Y(net67));
 INVx1_ASAP7_75t_SL _33 (.A(clknet_2_2__leaf_clock),
    .Y(net68));
 INVx1_ASAP7_75t_SL _33_34 (.A(clknet_2_2__leaf_clock),
    .Y(net69));
 INVx1_ASAP7_75t_SL _33_35 (.A(clknet_2_2__leaf_clock),
    .Y(net70));
 INVx1_ASAP7_75t_SL _33_36 (.A(clknet_2_2__leaf_clock),
    .Y(net71));
 INVx1_ASAP7_75t_SL _33_37 (.A(clknet_2_0__leaf_clock),
    .Y(net72));
 BUFx4_ASAP7_75t_SL clkbuf_2_0__f_clock (.A(clknet_0_clock),
    .Y(clknet_2_0__leaf_clock));
 BUFx4_ASAP7_75t_SL clkbuf_2_1__f_clock (.A(clknet_0_clock),
    .Y(clknet_2_1__leaf_clock));
 BUFx4_ASAP7_75t_SL clkbuf_2_2__f_clock (.A(clknet_0_clock),
    .Y(clknet_2_2__leaf_clock));
 BUFx4_ASAP7_75t_SL clkbuf_2_3__f_clock (.A(clknet_0_clock),
    .Y(clknet_2_3__leaf_clock));
 BUFx2_ASAP7_75t_SL rebuffer38 (.A(_033_),
    .Y(net73));
 BUFx2_ASAP7_75t_SL rebuffer39 (.A(_068_),
    .Y(net74));
 BUFx2_ASAP7_75t_SL rebuffer40 (.A(_067_),
    .Y(net75));
 DECAPx10_ASAP7_75t_SL FILLER_0_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_0_112 ();
 DECAPx2_ASAP7_75t_SL FILLER_0_120 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_0_126 ();
 DECAPx1_ASAP7_75t_SL FILLER_0_134 ();
 FILLERxp5_ASAP7_75t_SL FILLER_0_138 ();
 DECAPx4_ASAP7_75t_SL FILLER_0_144 ();
 FILLER_ASAP7_75t_SL FILLER_0_154 ();
 DECAPx2_ASAP7_75t_SL FILLER_0_161 ();
 FILLERxp5_ASAP7_75t_SL FILLER_0_167 ();
 DECAPx1_ASAP7_75t_SL FILLER_0_173 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_182 ();
 DECAPx2_ASAP7_75t_SL FILLER_0_204 ();
 FILLER_ASAP7_75t_SL FILLER_0_215 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_244 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_266 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_288 ();
 DECAPx4_ASAP7_75t_SL FILLER_0_310 ();
 FILLER_ASAP7_75t_SL FILLER_0_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_156 ();
 DECAPx6_ASAP7_75t_SL FILLER_1_178 ();
 DECAPx1_ASAP7_75t_SL FILLER_1_192 ();
 FILLERxp5_ASAP7_75t_SL FILLER_1_196 ();
 DECAPx2_ASAP7_75t_SL FILLER_1_202 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_1_208 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_216 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_238 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_260 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_282 ();
 DECAPx6_ASAP7_75t_SL FILLER_1_304 ();
 DECAPx1_ASAP7_75t_SL FILLER_1_318 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_244 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_266 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_288 ();
 DECAPx4_ASAP7_75t_SL FILLER_2_310 ();
 FILLER_ASAP7_75t_SL FILLER_2_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_244 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_266 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_288 ();
 DECAPx4_ASAP7_75t_SL FILLER_3_310 ();
 FILLER_ASAP7_75t_SL FILLER_3_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_244 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_266 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_288 ();
 DECAPx4_ASAP7_75t_SL FILLER_4_310 ();
 FILLER_ASAP7_75t_SL FILLER_4_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_244 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_266 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_288 ();
 DECAPx4_ASAP7_75t_SL FILLER_5_310 ();
 FILLER_ASAP7_75t_SL FILLER_5_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_112 ();
 DECAPx6_ASAP7_75t_SL FILLER_6_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_151 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_173 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_195 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_217 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_239 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_261 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_283 ();
 DECAPx6_ASAP7_75t_SL FILLER_6_305 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_6_319 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_90 ();
 DECAPx1_ASAP7_75t_SL FILLER_7_112 ();
 FILLERxp5_ASAP7_75t_SL FILLER_7_116 ();
 FILLER_ASAP7_75t_SL FILLER_7_138 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_161 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_183 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_205 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_227 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_249 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_271 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_293 ();
 DECAPx2_ASAP7_75t_SL FILLER_7_315 ();
 FILLERxp5_ASAP7_75t_SL FILLER_7_321 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_90 ();
 DECAPx6_ASAP7_75t_SL FILLER_8_112 ();
 FILLER_ASAP7_75t_SL FILLER_8_129 ();
 FILLER_ASAP7_75t_SL FILLER_8_137 ();
 DECAPx1_ASAP7_75t_SL FILLER_8_142 ();
 FILLERxp5_ASAP7_75t_SL FILLER_8_146 ();
 DECAPx2_ASAP7_75t_SL FILLER_8_153 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_162 ();
 DECAPx4_ASAP7_75t_SL FILLER_8_184 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_8_194 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_244 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_266 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_288 ();
 DECAPx4_ASAP7_75t_SL FILLER_8_310 ();
 FILLER_ASAP7_75t_SL FILLER_8_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_178 ();
 DECAPx1_ASAP7_75t_SL FILLER_9_200 ();
 FILLER_ASAP7_75t_SL FILLER_9_210 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_215 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_237 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_259 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_281 ();
 DECAPx6_ASAP7_75t_SL FILLER_9_303 ();
 DECAPx1_ASAP7_75t_SL FILLER_9_317 ();
 FILLERxp5_ASAP7_75t_SL FILLER_9_321 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_90 ();
 DECAPx4_ASAP7_75t_SL FILLER_10_112 ();
 FILLERxp5_ASAP7_75t_SL FILLER_10_122 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_126 ();
 DECAPx4_ASAP7_75t_SL FILLER_10_148 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_10_158 ();
 DECAPx6_ASAP7_75t_SL FILLER_10_164 ();
 FILLER_ASAP7_75t_SL FILLER_10_178 ();
 FILLER_ASAP7_75t_SL FILLER_10_201 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_224 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_246 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_268 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_290 ();
 DECAPx4_ASAP7_75t_SL FILLER_10_312 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_68 ();
 DECAPx6_ASAP7_75t_SL FILLER_11_90 ();
 FILLER_ASAP7_75t_SL FILLER_11_104 ();
 FILLER_ASAP7_75t_SL FILLER_11_127 ();
 DECAPx6_ASAP7_75t_SL FILLER_11_135 ();
 DECAPx1_ASAP7_75t_SL FILLER_11_149 ();
 DECAPx2_ASAP7_75t_SL FILLER_11_174 ();
 FILLER_ASAP7_75t_SL FILLER_11_180 ();
 DECAPx4_ASAP7_75t_SL FILLER_11_185 ();
 FILLER_ASAP7_75t_SL FILLER_11_195 ();
 FILLER_ASAP7_75t_SL FILLER_11_203 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_208 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_230 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_252 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_274 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_296 ();
 DECAPx1_ASAP7_75t_SL FILLER_11_318 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_68 ();
 DECAPx6_ASAP7_75t_SL FILLER_12_90 ();
 DECAPx1_ASAP7_75t_SL FILLER_12_104 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_111 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_133 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_158 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_180 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_12_202 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_226 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_248 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_270 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_292 ();
 DECAPx2_ASAP7_75t_SL FILLER_12_314 ();
 FILLER_ASAP7_75t_SL FILLER_12_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_134 ();
 DECAPx1_ASAP7_75t_SL FILLER_13_162 ();
 FILLER_ASAP7_75t_SL FILLER_13_172 ();
 DECAPx6_ASAP7_75t_SL FILLER_13_177 ();
 DECAPx1_ASAP7_75t_SL FILLER_13_191 ();
 FILLERxp5_ASAP7_75t_SL FILLER_13_195 ();
 DECAPx2_ASAP7_75t_SL FILLER_13_202 ();
 FILLER_ASAP7_75t_SL FILLER_13_214 ();
 FILLER_ASAP7_75t_SL FILLER_13_219 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_13_224 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_230 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_252 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_274 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_296 ();
 DECAPx1_ASAP7_75t_SL FILLER_13_318 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_112 ();
 DECAPx2_ASAP7_75t_SL FILLER_14_134 ();
 FILLER_ASAP7_75t_SL FILLER_14_140 ();
 FILLER_ASAP7_75t_SL FILLER_14_148 ();
 FILLER_ASAP7_75t_SL FILLER_14_156 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_14_179 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_14_188 ();
 DECAPx6_ASAP7_75t_SL FILLER_14_194 ();
 DECAPx1_ASAP7_75t_SL FILLER_14_208 ();
 FILLERxp5_ASAP7_75t_SL FILLER_14_212 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_234 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_256 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_278 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_300 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_134 ();
 DECAPx1_ASAP7_75t_SL FILLER_15_156 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_15_163 ();
 DECAPx1_ASAP7_75t_SL FILLER_15_173 ();
 DECAPx1_ASAP7_75t_SL FILLER_15_198 ();
 FILLER_ASAP7_75t_SL FILLER_15_208 ();
 FILLER_ASAP7_75t_SL FILLER_15_216 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_221 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_243 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_265 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_287 ();
 DECAPx4_ASAP7_75t_SL FILLER_15_309 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_15_319 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_134 ();
 DECAPx4_ASAP7_75t_SL FILLER_16_156 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_16_166 ();
 DECAPx1_ASAP7_75t_SL FILLER_16_175 ();
 DECAPx1_ASAP7_75t_SL FILLER_16_182 ();
 DECAPx4_ASAP7_75t_SL FILLER_16_192 ();
 FILLERxp5_ASAP7_75t_SL FILLER_16_202 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_209 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_231 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_253 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_275 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_297 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_16_319 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_134 ();
 DECAPx2_ASAP7_75t_SL FILLER_17_156 ();
 DECAPx6_ASAP7_75t_SL FILLER_17_168 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_17_182 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_244 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_266 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_288 ();
 DECAPx4_ASAP7_75t_SL FILLER_17_310 ();
 FILLER_ASAP7_75t_SL FILLER_17_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_18_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_18_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_18_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_18_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_18_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_18_112 ();
 DECAPx6_ASAP7_75t_SL FILLER_18_134 ();
 DECAPx1_ASAP7_75t_SL FILLER_18_148 ();
 DECAPx4_ASAP7_75t_SL FILLER_18_167 ();
 DECAPx2_ASAP7_75t_SL FILLER_18_183 ();
 FILLER_ASAP7_75t_SL FILLER_18_189 ();
 DECAPx6_ASAP7_75t_SL FILLER_18_206 ();
 FILLER_ASAP7_75t_SL FILLER_18_220 ();
 DECAPx10_ASAP7_75t_SL FILLER_18_229 ();
 DECAPx10_ASAP7_75t_SL FILLER_18_251 ();
 DECAPx10_ASAP7_75t_SL FILLER_18_273 ();
 DECAPx10_ASAP7_75t_SL FILLER_18_295 ();
 DECAPx1_ASAP7_75t_SL FILLER_18_317 ();
 FILLERxp5_ASAP7_75t_SL FILLER_18_321 ();
 DECAPx10_ASAP7_75t_SL FILLER_19_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_19_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_19_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_19_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_19_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_19_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_19_134 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_19_156 ();
 DECAPx6_ASAP7_75t_SL FILLER_19_174 ();
 DECAPx10_ASAP7_75t_SL FILLER_19_203 ();
 DECAPx10_ASAP7_75t_SL FILLER_19_225 ();
 DECAPx10_ASAP7_75t_SL FILLER_19_247 ();
 DECAPx10_ASAP7_75t_SL FILLER_19_269 ();
 DECAPx10_ASAP7_75t_SL FILLER_19_291 ();
 DECAPx2_ASAP7_75t_SL FILLER_19_313 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_19_319 ();
 DECAPx10_ASAP7_75t_SL FILLER_20_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_20_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_20_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_20_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_20_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_20_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_20_134 ();
 DECAPx6_ASAP7_75t_SL FILLER_20_156 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_20_170 ();
 FILLER_ASAP7_75t_SL FILLER_20_188 ();
 DECAPx4_ASAP7_75t_SL FILLER_20_196 ();
 FILLER_ASAP7_75t_SL FILLER_20_206 ();
 DECAPx10_ASAP7_75t_SL FILLER_20_214 ();
 DECAPx10_ASAP7_75t_SL FILLER_20_236 ();
 DECAPx10_ASAP7_75t_SL FILLER_20_258 ();
 DECAPx10_ASAP7_75t_SL FILLER_20_280 ();
 DECAPx6_ASAP7_75t_SL FILLER_20_302 ();
 DECAPx2_ASAP7_75t_SL FILLER_20_316 ();
 DECAPx10_ASAP7_75t_SL FILLER_21_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_21_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_21_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_21_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_21_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_21_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_21_134 ();
 DECAPx1_ASAP7_75t_SL FILLER_21_156 ();
 DECAPx6_ASAP7_75t_SL FILLER_21_175 ();
 DECAPx1_ASAP7_75t_SL FILLER_21_189 ();
 FILLERxp5_ASAP7_75t_SL FILLER_21_193 ();
 DECAPx10_ASAP7_75t_SL FILLER_21_209 ();
 DECAPx10_ASAP7_75t_SL FILLER_21_231 ();
 DECAPx6_ASAP7_75t_SL FILLER_21_253 ();
 DECAPx1_ASAP7_75t_SL FILLER_21_267 ();
 FILLERxp5_ASAP7_75t_SL FILLER_21_271 ();
 DECAPx10_ASAP7_75t_SL FILLER_21_293 ();
 DECAPx2_ASAP7_75t_SL FILLER_21_315 ();
 FILLERxp5_ASAP7_75t_SL FILLER_21_321 ();
 DECAPx2_ASAP7_75t_SL FILLER_22_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_22_8 ();
 DECAPx2_ASAP7_75t_SL FILLER_22_16 ();
 FILLERxp5_ASAP7_75t_SL FILLER_22_22 ();
 DECAPx10_ASAP7_75t_SL FILLER_22_28 ();
 DECAPx10_ASAP7_75t_SL FILLER_22_50 ();
 DECAPx10_ASAP7_75t_SL FILLER_22_72 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_22_94 ();
 DECAPx1_ASAP7_75t_SL FILLER_22_100 ();
 DECAPx10_ASAP7_75t_SL FILLER_22_125 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_22_147 ();
 FILLER_ASAP7_75t_SL FILLER_22_165 ();
 DECAPx6_ASAP7_75t_SL FILLER_22_173 ();
 DECAPx1_ASAP7_75t_SL FILLER_22_187 ();
 FILLERxp5_ASAP7_75t_SL FILLER_22_191 ();
 DECAPx10_ASAP7_75t_SL FILLER_22_198 ();
 DECAPx10_ASAP7_75t_SL FILLER_22_220 ();
 DECAPx10_ASAP7_75t_SL FILLER_22_242 ();
 DECAPx2_ASAP7_75t_SL FILLER_22_264 ();
 FILLER_ASAP7_75t_SL FILLER_22_270 ();
 FILLER_ASAP7_75t_SL FILLER_22_278 ();
 DECAPx2_ASAP7_75t_SL FILLER_22_283 ();
 DECAPx10_ASAP7_75t_SL FILLER_22_292 ();
 DECAPx2_ASAP7_75t_SL FILLER_22_314 ();
 FILLER_ASAP7_75t_SL FILLER_22_320 ();
 FILLER_ASAP7_75t_SL FILLER_23_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_23_9 ();
 DECAPx10_ASAP7_75t_SL FILLER_23_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_23_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_23_68 ();
 DECAPx6_ASAP7_75t_SL FILLER_23_90 ();
 FILLERxp5_ASAP7_75t_SL FILLER_23_104 ();
 DECAPx4_ASAP7_75t_SL FILLER_23_111 ();
 FILLER_ASAP7_75t_SL FILLER_23_121 ();
 DECAPx10_ASAP7_75t_SL FILLER_23_126 ();
 DECAPx6_ASAP7_75t_SL FILLER_23_148 ();
 DECAPx2_ASAP7_75t_SL FILLER_23_162 ();
 DECAPx2_ASAP7_75t_SL FILLER_23_183 ();
 DECAPx10_ASAP7_75t_SL FILLER_23_195 ();
 DECAPx10_ASAP7_75t_SL FILLER_23_217 ();
 DECAPx2_ASAP7_75t_SL FILLER_23_239 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_23_245 ();
 DECAPx10_ASAP7_75t_SL FILLER_23_254 ();
 DECAPx6_ASAP7_75t_SL FILLER_23_276 ();
 FILLERxp5_ASAP7_75t_SL FILLER_23_290 ();
 DECAPx10_ASAP7_75t_SL FILLER_23_296 ();
 DECAPx1_ASAP7_75t_SL FILLER_23_318 ();
 DECAPx10_ASAP7_75t_SL FILLER_24_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_24_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_24_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_24_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_24_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_24_112 ();
 DECAPx4_ASAP7_75t_SL FILLER_24_134 ();
 DECAPx4_ASAP7_75t_SL FILLER_24_150 ();
 FILLER_ASAP7_75t_SL FILLER_24_160 ();
 FILLER_ASAP7_75t_SL FILLER_24_168 ();
 DECAPx2_ASAP7_75t_SL FILLER_24_176 ();
 FILLER_ASAP7_75t_SL FILLER_24_182 ();
 DECAPx6_ASAP7_75t_SL FILLER_24_190 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_24_204 ();
 DECAPx6_ASAP7_75t_SL FILLER_24_213 ();
 FILLERxp5_ASAP7_75t_SL FILLER_24_227 ();
 DECAPx10_ASAP7_75t_SL FILLER_24_243 ();
 DECAPx10_ASAP7_75t_SL FILLER_24_265 ();
 DECAPx10_ASAP7_75t_SL FILLER_24_287 ();
 DECAPx4_ASAP7_75t_SL FILLER_24_309 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_24_319 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_112 ();
 DECAPx4_ASAP7_75t_SL FILLER_25_134 ();
 FILLER_ASAP7_75t_SL FILLER_25_159 ();
 DECAPx1_ASAP7_75t_SL FILLER_25_167 ();
 FILLERxp5_ASAP7_75t_SL FILLER_25_171 ();
 FILLER_ASAP7_75t_SL FILLER_25_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_186 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_208 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_230 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_252 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_274 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_296 ();
 DECAPx1_ASAP7_75t_SL FILLER_25_318 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_134 ();
 DECAPx2_ASAP7_75t_SL FILLER_26_156 ();
 FILLER_ASAP7_75t_SL FILLER_26_162 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_170 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_192 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_214 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_236 ();
 DECAPx4_ASAP7_75t_SL FILLER_26_258 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_26_268 ();
 DECAPx4_ASAP7_75t_SL FILLER_26_277 ();
 DECAPx4_ASAP7_75t_SL FILLER_26_290 ();
 FILLERxp5_ASAP7_75t_SL FILLER_26_300 ();
 DECAPx6_ASAP7_75t_SL FILLER_26_306 ();
 FILLER_ASAP7_75t_SL FILLER_26_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_90 ();
 DECAPx6_ASAP7_75t_SL FILLER_27_112 ();
 FILLERxp5_ASAP7_75t_SL FILLER_27_126 ();
 DECAPx6_ASAP7_75t_SL FILLER_27_142 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_27_156 ();
 FILLER_ASAP7_75t_SL FILLER_27_166 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_174 ();
 DECAPx6_ASAP7_75t_SL FILLER_27_196 ();
 DECAPx1_ASAP7_75t_SL FILLER_27_210 ();
 FILLER_ASAP7_75t_SL FILLER_27_220 ();
 DECAPx2_ASAP7_75t_SL FILLER_27_237 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_27_243 ();
 DECAPx6_ASAP7_75t_SL FILLER_27_252 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_27_266 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_290 ();
 DECAPx4_ASAP7_75t_SL FILLER_27_312 ();
 DECAPx10_ASAP7_75t_SL FILLER_28_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_28_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_28_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_28_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_28_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_28_112 ();
 DECAPx2_ASAP7_75t_SL FILLER_28_134 ();
 FILLERxp5_ASAP7_75t_SL FILLER_28_140 ();
 DECAPx2_ASAP7_75t_SL FILLER_28_147 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_28_153 ();
 FILLER_ASAP7_75t_SL FILLER_28_168 ();
 DECAPx1_ASAP7_75t_SL FILLER_28_177 ();
 DECAPx6_ASAP7_75t_SL FILLER_28_188 ();
 DECAPx2_ASAP7_75t_SL FILLER_28_202 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_28_214 ();
 DECAPx1_ASAP7_75t_SL FILLER_28_223 ();
 FILLERxp5_ASAP7_75t_SL FILLER_28_227 ();
 DECAPx2_ASAP7_75t_SL FILLER_28_243 ();
 FILLERxp5_ASAP7_75t_SL FILLER_28_249 ();
 DECAPx4_ASAP7_75t_SL FILLER_28_256 ();
 FILLER_ASAP7_75t_SL FILLER_28_272 ();
 DECAPx2_ASAP7_75t_SL FILLER_28_277 ();
 FILLER_ASAP7_75t_SL FILLER_28_286 ();
 DECAPx4_ASAP7_75t_SL FILLER_28_294 ();
 FILLER_ASAP7_75t_SL FILLER_28_304 ();
 FILLER_ASAP7_75t_SL FILLER_28_311 ();
 DECAPx1_ASAP7_75t_SL FILLER_28_318 ();
 DECAPx10_ASAP7_75t_SL FILLER_29_2 ();
 FILLER_ASAP7_75t_SL FILLER_29_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_29_31 ();
 DECAPx10_ASAP7_75t_SL FILLER_29_53 ();
 DECAPx10_ASAP7_75t_SL FILLER_29_75 ();
 DECAPx10_ASAP7_75t_SL FILLER_29_97 ();
 DECAPx1_ASAP7_75t_SL FILLER_29_119 ();
 DECAPx1_ASAP7_75t_SL FILLER_29_129 ();
 FILLERxp5_ASAP7_75t_SL FILLER_29_133 ();
 DECAPx10_ASAP7_75t_SL FILLER_29_137 ();
 FILLER_ASAP7_75t_SL FILLER_29_179 ();
 DECAPx10_ASAP7_75t_SL FILLER_29_187 ();
 DECAPx6_ASAP7_75t_SL FILLER_29_209 ();
 DECAPx1_ASAP7_75t_SL FILLER_29_223 ();
 FILLER_ASAP7_75t_SL FILLER_29_242 ();
 DECAPx6_ASAP7_75t_SL FILLER_29_250 ();
 FILLER_ASAP7_75t_SL FILLER_29_264 ();
 FILLER_ASAP7_75t_SL FILLER_29_287 ();
 FILLER_ASAP7_75t_SL FILLER_29_310 ();
 DECAPx2_ASAP7_75t_SL FILLER_29_315 ();
 FILLERxp5_ASAP7_75t_SL FILLER_29_321 ();
 DECAPx10_ASAP7_75t_SL FILLER_30_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_30_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_30_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_30_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_30_90 ();
 DECAPx1_ASAP7_75t_SL FILLER_30_112 ();
 FILLERxp5_ASAP7_75t_SL FILLER_30_116 ();
 DECAPx6_ASAP7_75t_SL FILLER_30_138 ();
 FILLERxp5_ASAP7_75t_SL FILLER_30_152 ();
 FILLER_ASAP7_75t_SL FILLER_30_159 ();
 FILLER_ASAP7_75t_SL FILLER_30_167 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_30_176 ();
 FILLER_ASAP7_75t_SL FILLER_30_184 ();
 FILLER_ASAP7_75t_SL FILLER_30_193 ();
 DECAPx10_ASAP7_75t_SL FILLER_30_198 ();
 DECAPx10_ASAP7_75t_SL FILLER_30_220 ();
 DECAPx10_ASAP7_75t_SL FILLER_30_242 ();
 DECAPx1_ASAP7_75t_SL FILLER_30_264 ();
 DECAPx6_ASAP7_75t_SL FILLER_30_271 ();
 DECAPx2_ASAP7_75t_SL FILLER_30_285 ();
 DECAPx10_ASAP7_75t_SL FILLER_30_294 ();
 DECAPx2_ASAP7_75t_SL FILLER_30_316 ();
 DECAPx10_ASAP7_75t_SL FILLER_31_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_31_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_31_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_31_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_31_90 ();
 DECAPx2_ASAP7_75t_SL FILLER_31_112 ();
 FILLERxp5_ASAP7_75t_SL FILLER_31_118 ();
 DECAPx10_ASAP7_75t_SL FILLER_31_122 ();
 DECAPx4_ASAP7_75t_SL FILLER_31_144 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_31_160 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_31_166 ();
 FILLER_ASAP7_75t_SL FILLER_31_172 ();
 FILLER_ASAP7_75t_SL FILLER_31_189 ();
 DECAPx4_ASAP7_75t_SL FILLER_31_206 ();
 FILLER_ASAP7_75t_SL FILLER_31_222 ();
 DECAPx1_ASAP7_75t_SL FILLER_31_239 ();
 DECAPx10_ASAP7_75t_SL FILLER_31_249 ();
 DECAPx10_ASAP7_75t_SL FILLER_31_271 ();
 DECAPx10_ASAP7_75t_SL FILLER_31_293 ();
 DECAPx2_ASAP7_75t_SL FILLER_31_315 ();
 FILLERxp5_ASAP7_75t_SL FILLER_31_321 ();
 DECAPx10_ASAP7_75t_SL FILLER_32_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_32_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_32_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_32_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_32_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_32_112 ();
 DECAPx4_ASAP7_75t_SL FILLER_32_134 ();
 FILLERxp5_ASAP7_75t_SL FILLER_32_144 ();
 DECAPx1_ASAP7_75t_SL FILLER_32_165 ();
 FILLER_ASAP7_75t_SL FILLER_32_176 ();
 DECAPx2_ASAP7_75t_SL FILLER_32_183 ();
 FILLER_ASAP7_75t_SL FILLER_32_195 ();
 DECAPx2_ASAP7_75t_SL FILLER_32_201 ();
 FILLERxp5_ASAP7_75t_SL FILLER_32_207 ();
 FILLER_ASAP7_75t_SL FILLER_32_214 ();
 DECAPx10_ASAP7_75t_SL FILLER_32_222 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_32_244 ();
 DECAPx2_ASAP7_75t_SL FILLER_32_253 ();
 FILLER_ASAP7_75t_SL FILLER_32_265 ();
 FILLER_ASAP7_75t_SL FILLER_32_288 ();
 DECAPx2_ASAP7_75t_SL FILLER_32_293 ();
 FILLER_ASAP7_75t_SL FILLER_32_299 ();
 FILLER_ASAP7_75t_SL FILLER_32_306 ();
 DECAPx2_ASAP7_75t_SL FILLER_32_313 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_32_319 ();
 DECAPx10_ASAP7_75t_SL FILLER_33_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_33_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_33_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_33_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_33_90 ();
 DECAPx4_ASAP7_75t_SL FILLER_33_112 ();
 FILLER_ASAP7_75t_SL FILLER_33_122 ();
 FILLER_ASAP7_75t_SL FILLER_33_145 ();
 DECAPx1_ASAP7_75t_SL FILLER_33_150 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_33_174 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_33_183 ();
 DECAPx6_ASAP7_75t_SL FILLER_33_195 ();
 DECAPx1_ASAP7_75t_SL FILLER_33_215 ();
 FILLERxp5_ASAP7_75t_SL FILLER_33_219 ();
 FILLER_ASAP7_75t_SL FILLER_33_235 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_33_243 ();
 FILLER_ASAP7_75t_SL FILLER_33_267 ();
 DECAPx1_ASAP7_75t_SL FILLER_33_272 ();
 DECAPx10_ASAP7_75t_SL FILLER_33_282 ();
 DECAPx6_ASAP7_75t_SL FILLER_33_304 ();
 DECAPx1_ASAP7_75t_SL FILLER_33_318 ();
 DECAPx4_ASAP7_75t_SL FILLER_34_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_34_12 ();
 DECAPx10_ASAP7_75t_SL FILLER_34_20 ();
 DECAPx10_ASAP7_75t_SL FILLER_34_42 ();
 DECAPx10_ASAP7_75t_SL FILLER_34_64 ();
 DECAPx6_ASAP7_75t_SL FILLER_34_86 ();
 DECAPx2_ASAP7_75t_SL FILLER_34_100 ();
 FILLERxp5_ASAP7_75t_SL FILLER_34_106 ();
 FILLER_ASAP7_75t_SL FILLER_34_113 ();
 DECAPx2_ASAP7_75t_SL FILLER_34_118 ();
 FILLERxp5_ASAP7_75t_SL FILLER_34_124 ();
 FILLER_ASAP7_75t_SL FILLER_34_128 ();
 DECAPx1_ASAP7_75t_SL FILLER_34_136 ();
 FILLERxp5_ASAP7_75t_SL FILLER_34_140 ();
 FILLER_ASAP7_75t_SL FILLER_34_144 ();
 FILLER_ASAP7_75t_SL FILLER_34_152 ();
 FILLER_ASAP7_75t_SL FILLER_34_160 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_34_168 ();
 FILLER_ASAP7_75t_SL FILLER_34_176 ();
 FILLER_ASAP7_75t_SL FILLER_34_184 ();
 DECAPx2_ASAP7_75t_SL FILLER_34_189 ();
 FILLER_ASAP7_75t_SL FILLER_34_195 ();
 FILLER_ASAP7_75t_SL FILLER_34_204 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_34_212 ();
 FILLER_ASAP7_75t_SL FILLER_34_221 ();
 DECAPx4_ASAP7_75t_SL FILLER_34_238 ();
 DECAPx6_ASAP7_75t_SL FILLER_34_251 ();
 DECAPx1_ASAP7_75t_SL FILLER_34_265 ();
 DECAPx1_ASAP7_75t_SL FILLER_34_272 ();
 FILLER_ASAP7_75t_SL FILLER_34_297 ();
 DECAPx6_ASAP7_75t_SL FILLER_34_302 ();
 DECAPx2_ASAP7_75t_SL FILLER_34_316 ();
 DECAPx4_ASAP7_75t_SL FILLER_35_2 ();
 FILLERxp5_ASAP7_75t_SL FILLER_35_12 ();
 DECAPx10_ASAP7_75t_SL FILLER_35_18 ();
 DECAPx10_ASAP7_75t_SL FILLER_35_40 ();
 DECAPx10_ASAP7_75t_SL FILLER_35_62 ();
 DECAPx6_ASAP7_75t_SL FILLER_35_84 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_35_98 ();
 DECAPx10_ASAP7_75t_SL FILLER_35_122 ();
 DECAPx6_ASAP7_75t_SL FILLER_35_144 ();
 FILLERxp5_ASAP7_75t_SL FILLER_35_158 ();
 FILLER_ASAP7_75t_SL FILLER_35_174 ();
 DECAPx10_ASAP7_75t_SL FILLER_35_186 ();
 DECAPx6_ASAP7_75t_SL FILLER_35_208 ();
 FILLER_ASAP7_75t_SL FILLER_35_222 ();
 DECAPx4_ASAP7_75t_SL FILLER_35_239 ();
 DECAPx6_ASAP7_75t_SL FILLER_35_255 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_35_269 ();
 FILLER_ASAP7_75t_SL FILLER_35_275 ();
 FILLER_ASAP7_75t_SL FILLER_35_298 ();
 FILLER_ASAP7_75t_SL FILLER_35_303 ();
 DECAPx4_ASAP7_75t_SL FILLER_35_310 ();
 FILLER_ASAP7_75t_SL FILLER_35_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_36_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_36_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_36_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_36_68 ();
 DECAPx4_ASAP7_75t_SL FILLER_36_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_36_100 ();
 DECAPx10_ASAP7_75t_SL FILLER_36_106 ();
 DECAPx10_ASAP7_75t_SL FILLER_36_128 ();
 DECAPx2_ASAP7_75t_SL FILLER_36_150 ();
 FILLER_ASAP7_75t_SL FILLER_36_156 ();
 DECAPx4_ASAP7_75t_SL FILLER_36_168 ();
 FILLER_ASAP7_75t_SL FILLER_36_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_36_190 ();
 DECAPx1_ASAP7_75t_SL FILLER_36_212 ();
 FILLERxp5_ASAP7_75t_SL FILLER_36_216 ();
 DECAPx6_ASAP7_75t_SL FILLER_36_232 ();
 FILLERxp5_ASAP7_75t_SL FILLER_36_246 ();
 DECAPx4_ASAP7_75t_SL FILLER_36_253 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_36_263 ();
 FILLER_ASAP7_75t_SL FILLER_36_272 ();
 FILLER_ASAP7_75t_SL FILLER_36_295 ();
 DECAPx2_ASAP7_75t_SL FILLER_36_300 ();
 FILLER_ASAP7_75t_SL FILLER_36_306 ();
 DECAPx2_ASAP7_75t_SL FILLER_36_313 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_36_319 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_222 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_37_244 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_253 ();
 FILLER_ASAP7_75t_SL FILLER_37_275 ();
 FILLER_ASAP7_75t_SL FILLER_37_283 ();
 DECAPx1_ASAP7_75t_SL FILLER_37_288 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_295 ();
 DECAPx1_ASAP7_75t_SL FILLER_37_317 ();
 FILLERxp5_ASAP7_75t_SL FILLER_37_321 ();
 DECAPx10_ASAP7_75t_SL FILLER_38_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_38_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_38_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_38_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_38_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_38_112 ();
 DECAPx2_ASAP7_75t_SL FILLER_38_134 ();
 DECAPx6_ASAP7_75t_SL FILLER_38_152 ();
 FILLERxp5_ASAP7_75t_SL FILLER_38_166 ();
 DECAPx10_ASAP7_75t_SL FILLER_38_177 ();
 DECAPx6_ASAP7_75t_SL FILLER_38_199 ();
 DECAPx1_ASAP7_75t_SL FILLER_38_213 ();
 DECAPx6_ASAP7_75t_SL FILLER_38_255 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_38_269 ();
 DECAPx10_ASAP7_75t_SL FILLER_38_278 ();
 DECAPx6_ASAP7_75t_SL FILLER_38_305 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_38_319 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_112 ();
 DECAPx4_ASAP7_75t_SL FILLER_39_134 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_39_144 ();
 DECAPx4_ASAP7_75t_SL FILLER_39_153 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_39_163 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_170 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_192 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_214 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_236 ();
 DECAPx6_ASAP7_75t_SL FILLER_39_258 ();
 FILLER_ASAP7_75t_SL FILLER_39_293 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_298 ();
 FILLER_ASAP7_75t_SL FILLER_39_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_112 ();
 DECAPx4_ASAP7_75t_SL FILLER_40_134 ();
 FILLER_ASAP7_75t_SL FILLER_40_144 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_166 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_188 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_210 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_232 ();
 DECAPx6_ASAP7_75t_SL FILLER_40_254 ();
 DECAPx2_ASAP7_75t_SL FILLER_40_268 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_277 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_299 ();
 FILLERxp5_ASAP7_75t_SL FILLER_40_321 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_112 ();
 DECAPx6_ASAP7_75t_SL FILLER_41_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_151 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_173 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_195 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_217 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_239 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_261 ();
 DECAPx6_ASAP7_75t_SL FILLER_41_283 ();
 DECAPx1_ASAP7_75t_SL FILLER_41_297 ();
 DECAPx6_ASAP7_75t_SL FILLER_41_306 ();
 FILLER_ASAP7_75t_SL FILLER_41_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_112 ();
 DECAPx6_ASAP7_75t_SL FILLER_42_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_154 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_176 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_198 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_220 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_242 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_264 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_286 ();
 DECAPx6_ASAP7_75t_SL FILLER_42_308 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_112 ();
 DECAPx6_ASAP7_75t_SL FILLER_43_134 ();
 FILLER_ASAP7_75t_SL FILLER_43_155 ();
 FILLER_ASAP7_75t_SL FILLER_43_163 ();
 DECAPx2_ASAP7_75t_SL FILLER_43_171 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_43_177 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_186 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_208 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_230 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_252 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_274 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_296 ();
 DECAPx1_ASAP7_75t_SL FILLER_43_318 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_112 ();
 DECAPx2_ASAP7_75t_SL FILLER_44_134 ();
 FILLERxp5_ASAP7_75t_SL FILLER_44_140 ();
 FILLER_ASAP7_75t_SL FILLER_44_147 ();
 FILLER_ASAP7_75t_SL FILLER_44_164 ();
 DECAPx2_ASAP7_75t_SL FILLER_44_172 ();
 FILLERxp5_ASAP7_75t_SL FILLER_44_178 ();
 DECAPx6_ASAP7_75t_SL FILLER_44_182 ();
 DECAPx2_ASAP7_75t_SL FILLER_44_196 ();
 FILLERxp5_ASAP7_75t_SL FILLER_44_202 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_210 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_232 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_254 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_276 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_298 ();
 FILLER_ASAP7_75t_SL FILLER_44_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_112 ();
 FILLER_ASAP7_75t_SL FILLER_45_134 ();
 FILLER_ASAP7_75t_SL FILLER_45_142 ();
 FILLER_ASAP7_75t_SL FILLER_45_152 ();
 FILLER_ASAP7_75t_SL FILLER_45_160 ();
 DECAPx2_ASAP7_75t_SL FILLER_45_168 ();
 FILLER_ASAP7_75t_SL FILLER_45_174 ();
 FILLER_ASAP7_75t_SL FILLER_45_182 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_199 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_221 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_243 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_265 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_287 ();
 DECAPx4_ASAP7_75t_SL FILLER_45_309 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_45_319 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_90 ();
 DECAPx6_ASAP7_75t_SL FILLER_46_112 ();
 FILLERxp5_ASAP7_75t_SL FILLER_46_126 ();
 DECAPx1_ASAP7_75t_SL FILLER_46_147 ();
 DECAPx2_ASAP7_75t_SL FILLER_46_166 ();
 FILLERxp5_ASAP7_75t_SL FILLER_46_172 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_188 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_210 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_232 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_254 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_276 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_298 ();
 FILLER_ASAP7_75t_SL FILLER_46_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_90 ();
 DECAPx6_ASAP7_75t_SL FILLER_47_112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_47_126 ();
 DECAPx6_ASAP7_75t_SL FILLER_47_132 ();
 DECAPx2_ASAP7_75t_SL FILLER_47_161 ();
 FILLER_ASAP7_75t_SL FILLER_47_167 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_184 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_206 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_228 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_250 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_272 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_294 ();
 DECAPx2_ASAP7_75t_SL FILLER_47_316 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_112 ();
 DECAPx4_ASAP7_75t_SL FILLER_48_134 ();
 FILLER_ASAP7_75t_SL FILLER_48_159 ();
 FILLER_ASAP7_75t_SL FILLER_48_167 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_184 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_206 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_228 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_250 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_272 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_294 ();
 DECAPx2_ASAP7_75t_SL FILLER_48_316 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_112 ();
 DECAPx6_ASAP7_75t_SL FILLER_49_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_154 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_176 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_198 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_220 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_242 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_264 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_286 ();
 DECAPx6_ASAP7_75t_SL FILLER_49_308 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_134 ();
 FILLERxp5_ASAP7_75t_SL FILLER_50_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_163 ();
 FILLERxp5_ASAP7_75t_SL FILLER_50_185 ();
 DECAPx2_ASAP7_75t_SL FILLER_50_192 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_204 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_226 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_248 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_270 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_292 ();
 DECAPx2_ASAP7_75t_SL FILLER_50_314 ();
 FILLER_ASAP7_75t_SL FILLER_50_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_134 ();
 DECAPx1_ASAP7_75t_SL FILLER_51_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_166 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_188 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_210 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_232 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_254 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_276 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_298 ();
 FILLER_ASAP7_75t_SL FILLER_51_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_134 ();
 FILLER_ASAP7_75t_SL FILLER_52_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_164 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_186 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_208 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_230 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_252 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_274 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_296 ();
 DECAPx1_ASAP7_75t_SL FILLER_52_318 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_134 ();
 FILLER_ASAP7_75t_SL FILLER_53_156 ();
 DECAPx1_ASAP7_75t_SL FILLER_53_179 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_189 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_211 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_233 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_255 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_277 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_299 ();
 FILLERxp5_ASAP7_75t_SL FILLER_53_321 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_112 ();
 DECAPx2_ASAP7_75t_SL FILLER_54_134 ();
 FILLERxp5_ASAP7_75t_SL FILLER_54_140 ();
 FILLER_ASAP7_75t_SL FILLER_54_147 ();
 DECAPx1_ASAP7_75t_SL FILLER_54_152 ();
 FILLER_ASAP7_75t_SL FILLER_54_159 ();
 FILLER_ASAP7_75t_SL FILLER_54_167 ();
 DECAPx2_ASAP7_75t_SL FILLER_54_172 ();
 FILLER_ASAP7_75t_SL FILLER_54_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_186 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_208 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_230 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_252 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_274 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_296 ();
 DECAPx1_ASAP7_75t_SL FILLER_54_318 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_112 ();
 FILLERxp5_ASAP7_75t_SL FILLER_55_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_156 ();
 FILLERxp5_ASAP7_75t_SL FILLER_55_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_244 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_266 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_288 ();
 DECAPx4_ASAP7_75t_SL FILLER_55_310 ();
 FILLER_ASAP7_75t_SL FILLER_55_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_56_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_56_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_56_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_56_68 ();
 DECAPx6_ASAP7_75t_SL FILLER_56_90 ();
 DECAPx2_ASAP7_75t_SL FILLER_56_104 ();
 FILLERxp5_ASAP7_75t_SL FILLER_56_110 ();
 FILLER_ASAP7_75t_SL FILLER_56_132 ();
 FILLER_ASAP7_75t_SL FILLER_56_140 ();
 DECAPx10_ASAP7_75t_SL FILLER_56_145 ();
 DECAPx1_ASAP7_75t_SL FILLER_56_167 ();
 FILLERxp5_ASAP7_75t_SL FILLER_56_171 ();
 FILLER_ASAP7_75t_SL FILLER_56_175 ();
 FILLER_ASAP7_75t_SL FILLER_56_183 ();
 DECAPx10_ASAP7_75t_SL FILLER_56_206 ();
 DECAPx10_ASAP7_75t_SL FILLER_56_228 ();
 DECAPx10_ASAP7_75t_SL FILLER_56_250 ();
 DECAPx10_ASAP7_75t_SL FILLER_56_272 ();
 DECAPx10_ASAP7_75t_SL FILLER_56_294 ();
 DECAPx2_ASAP7_75t_SL FILLER_56_316 ();
 DECAPx10_ASAP7_75t_SL FILLER_57_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_57_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_57_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_57_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_57_90 ();
 FILLERxp5_ASAP7_75t_SL FILLER_57_112 ();
 DECAPx4_ASAP7_75t_SL FILLER_57_116 ();
 FILLER_ASAP7_75t_SL FILLER_57_126 ();
 DECAPx10_ASAP7_75t_SL FILLER_57_131 ();
 FILLER_ASAP7_75t_SL FILLER_57_153 ();
 DECAPx2_ASAP7_75t_SL FILLER_57_176 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_57_182 ();
 FILLER_ASAP7_75t_SL FILLER_57_191 ();
 FILLER_ASAP7_75t_SL FILLER_57_196 ();
 FILLER_ASAP7_75t_SL FILLER_57_201 ();
 DECAPx10_ASAP7_75t_SL FILLER_57_206 ();
 DECAPx10_ASAP7_75t_SL FILLER_57_228 ();
 DECAPx10_ASAP7_75t_SL FILLER_57_250 ();
 DECAPx10_ASAP7_75t_SL FILLER_57_272 ();
 DECAPx10_ASAP7_75t_SL FILLER_57_294 ();
 DECAPx2_ASAP7_75t_SL FILLER_57_316 ();
 DECAPx10_ASAP7_75t_SL FILLER_58_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_58_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_58_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_58_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_58_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_58_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_58_134 ();
 FILLERxp5_ASAP7_75t_SL FILLER_58_156 ();
 DECAPx1_ASAP7_75t_SL FILLER_58_160 ();
 FILLERxp5_ASAP7_75t_SL FILLER_58_164 ();
 FILLER_ASAP7_75t_SL FILLER_58_168 ();
 DECAPx1_ASAP7_75t_SL FILLER_58_191 ();
 FILLER_ASAP7_75t_SL FILLER_58_198 ();
 DECAPx10_ASAP7_75t_SL FILLER_58_206 ();
 DECAPx10_ASAP7_75t_SL FILLER_58_228 ();
 DECAPx10_ASAP7_75t_SL FILLER_58_250 ();
 DECAPx10_ASAP7_75t_SL FILLER_58_272 ();
 DECAPx10_ASAP7_75t_SL FILLER_58_294 ();
 DECAPx2_ASAP7_75t_SL FILLER_58_316 ();
 DECAPx10_ASAP7_75t_SL FILLER_59_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_59_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_59_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_59_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_59_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_59_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_59_134 ();
 DECAPx6_ASAP7_75t_SL FILLER_59_156 ();
 FILLER_ASAP7_75t_SL FILLER_59_170 ();
 DECAPx2_ASAP7_75t_SL FILLER_59_175 ();
 DECAPx6_ASAP7_75t_SL FILLER_59_187 ();
 DECAPx10_ASAP7_75t_SL FILLER_59_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_59_244 ();
 DECAPx10_ASAP7_75t_SL FILLER_59_266 ();
 DECAPx10_ASAP7_75t_SL FILLER_59_288 ();
 DECAPx4_ASAP7_75t_SL FILLER_59_310 ();
 FILLER_ASAP7_75t_SL FILLER_59_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_60_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_60_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_60_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_60_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_60_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_60_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_60_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_60_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_60_178 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_60_200 ();
 FILLER_ASAP7_75t_SL FILLER_60_206 ();
 DECAPx10_ASAP7_75t_SL FILLER_60_211 ();
 DECAPx10_ASAP7_75t_SL FILLER_60_233 ();
 DECAPx10_ASAP7_75t_SL FILLER_60_255 ();
 DECAPx10_ASAP7_75t_SL FILLER_60_277 ();
 DECAPx10_ASAP7_75t_SL FILLER_60_299 ();
 FILLERxp5_ASAP7_75t_SL FILLER_60_321 ();
 DECAPx10_ASAP7_75t_SL FILLER_61_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_61_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_61_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_61_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_61_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_61_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_61_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_61_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_61_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_61_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_61_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_61_244 ();
 DECAPx10_ASAP7_75t_SL FILLER_61_266 ();
 DECAPx10_ASAP7_75t_SL FILLER_61_288 ();
 DECAPx4_ASAP7_75t_SL FILLER_61_310 ();
 FILLER_ASAP7_75t_SL FILLER_61_320 ();
 DECAPx10_ASAP7_75t_SL FILLER_62_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_62_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_62_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_62_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_62_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_62_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_62_134 ();
 FILLERxp5_ASAP7_75t_SL FILLER_62_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_62_162 ();
 DECAPx1_ASAP7_75t_SL FILLER_62_184 ();
 FILLERxp5_ASAP7_75t_SL FILLER_62_188 ();
 FILLER_ASAP7_75t_SL FILLER_62_194 ();
 DECAPx2_ASAP7_75t_SL FILLER_62_201 ();
 FILLERxp5_ASAP7_75t_SL FILLER_62_207 ();
 DECAPx10_ASAP7_75t_SL FILLER_62_230 ();
 DECAPx10_ASAP7_75t_SL FILLER_62_252 ();
 DECAPx10_ASAP7_75t_SL FILLER_62_274 ();
 DECAPx10_ASAP7_75t_SL FILLER_62_296 ();
 DECAPx1_ASAP7_75t_SL FILLER_62_318 ();
 DECAPx10_ASAP7_75t_SL FILLER_63_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_63_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_63_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_63_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_63_90 ();
 DECAPx2_ASAP7_75t_SL FILLER_63_112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_63_118 ();
 DECAPx2_ASAP7_75t_SL FILLER_63_126 ();
 DECAPx10_ASAP7_75t_SL FILLER_63_137 ();
 FILLERxp5_ASAP7_75t_SL FILLER_63_159 ();
 DECAPx6_ASAP7_75t_SL FILLER_63_165 ();
 DECAPx6_ASAP7_75t_SL FILLER_63_184 ();
 FILLER_ASAP7_75t_SL FILLER_63_198 ();
 DECAPx10_ASAP7_75t_SL FILLER_63_205 ();
 DECAPx10_ASAP7_75t_SL FILLER_63_227 ();
 DECAPx10_ASAP7_75t_SL FILLER_63_249 ();
 DECAPx10_ASAP7_75t_SL FILLER_63_271 ();
 DECAPx10_ASAP7_75t_SL FILLER_63_293 ();
 DECAPx2_ASAP7_75t_SL FILLER_63_315 ();
 FILLERxp5_ASAP7_75t_SL FILLER_63_321 ();
endmodule
