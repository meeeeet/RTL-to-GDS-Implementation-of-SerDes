module ser (clock,
    dout,
    enable,
    load,
    din);
 input clock;
 output dout;
 input enable;
 input load;
 input [31:0] din;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire clknet_0_clock;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire net10;
 wire net9;
 wire _078_;
 wire net8;
 wire net7;
 wire net6;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire net5;
 wire net4;
 wire _139_;
 wire net3;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire net2;
 wire _149_;
 wire _150_;
 wire _151_;
 wire net1;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire clknet_2_0__leaf_clock;
 wire clknet_2_1__leaf_clock;
 wire clknet_2_2__leaf_clock;
 wire clknet_2_3__leaf_clock;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;

 INVx1_ASAP7_75t_SL _183_ (.A(net33),
    .Y(_075_));
 TAPCELL_ASAP7_75t_SL PHY_11 ();
 TAPCELL_ASAP7_75t_SL PHY_10 ();
 CKINVDCx6p67_ASAP7_75t_SL _186_ (.A(net74),
    .Y(_078_));
 TAPCELL_ASAP7_75t_SL PHY_9 ();
 TAPCELL_ASAP7_75t_SL PHY_8 ();
 TAPCELL_ASAP7_75t_SL PHY_7 ();
 AND2x2_ASAP7_75t_SL _190_ (.A(net73),
    .B(_009_),
    .Y(_082_));
 AO21x1_ASAP7_75t_SL _191_ (.A1(_078_),
    .A2(_008_),
    .B(_082_),
    .Y(_083_));
 AND3x1_ASAP7_75t_SL _192_ (.A(net76),
    .B(net78),
    .C(_083_),
    .Y(_084_));
 INVx1_ASAP7_75t_SL _193_ (.A(_000_),
    .Y(_085_));
 AND2x2_ASAP7_75t_SL _194_ (.A(_036_),
    .B(_085_),
    .Y(_086_));
 AND2x2_ASAP7_75t_SL _195_ (.A(net73),
    .B(_005_),
    .Y(_087_));
 AO21x1_ASAP7_75t_SL _196_ (.A1(_078_),
    .A2(_004_),
    .B(_087_),
    .Y(_088_));
 NOR2x1_ASAP7_75t_SL _197_ (.A(net77),
    .B(net78),
    .Y(_089_));
 AND2x2_ASAP7_75t_SL _198_ (.A(net73),
    .B(_003_),
    .Y(_090_));
 AO21x1_ASAP7_75t_SL _199_ (.A1(_078_),
    .A2(_002_),
    .B(_090_),
    .Y(_091_));
 AO22x1_ASAP7_75t_SL _200_ (.A1(_086_),
    .A2(_088_),
    .B1(_089_),
    .B2(_091_),
    .Y(_092_));
 INVx2_ASAP7_75t_SL _201_ (.A(net76),
    .Y(_093_));
 AND2x2_ASAP7_75t_SL _202_ (.A(net73),
    .B(_007_),
    .Y(_094_));
 AO21x1_ASAP7_75t_SL _203_ (.A1(_078_),
    .A2(_006_),
    .B(_094_),
    .Y(_095_));
 AND3x1_ASAP7_75t_SL _204_ (.A(_093_),
    .B(net78),
    .C(_095_),
    .Y(_096_));
 OR5x1_ASAP7_75t_SL _205_ (.A(_035_),
    .B(_034_),
    .C(_084_),
    .D(_092_),
    .E(_096_),
    .Y(_097_));
 INVx1_ASAP7_75t_SL _206_ (.A(_035_),
    .Y(_098_));
 AND2x2_ASAP7_75t_SL _207_ (.A(net73),
    .B(_017_),
    .Y(_099_));
 AO21x1_ASAP7_75t_SL _208_ (.A1(_078_),
    .A2(_016_),
    .B(_099_),
    .Y(_100_));
 AND3x1_ASAP7_75t_SL _209_ (.A(net76),
    .B(net78),
    .C(_100_),
    .Y(_101_));
 AND2x2_ASAP7_75t_SL _210_ (.A(net73),
    .B(_013_),
    .Y(_102_));
 AO21x1_ASAP7_75t_SL _211_ (.A1(_078_),
    .A2(_012_),
    .B(_102_),
    .Y(_103_));
 AND2x2_ASAP7_75t_SL _212_ (.A(net73),
    .B(_011_),
    .Y(_104_));
 AO21x1_ASAP7_75t_SL _213_ (.A1(_078_),
    .A2(_010_),
    .B(_104_),
    .Y(_105_));
 AO22x1_ASAP7_75t_SL _214_ (.A1(_086_),
    .A2(_103_),
    .B1(_105_),
    .B2(_089_),
    .Y(_106_));
 AND2x2_ASAP7_75t_SL _215_ (.A(net73),
    .B(_015_),
    .Y(_107_));
 AO21x1_ASAP7_75t_SL _216_ (.A1(_078_),
    .A2(_014_),
    .B(_107_),
    .Y(_108_));
 AND3x1_ASAP7_75t_SL _217_ (.A(_093_),
    .B(net78),
    .C(_108_),
    .Y(_109_));
 OR5x1_ASAP7_75t_SL _218_ (.A(_098_),
    .B(_034_),
    .C(_101_),
    .D(_106_),
    .E(_109_),
    .Y(_110_));
 INVx1_ASAP7_75t_SL _219_ (.A(_034_),
    .Y(_111_));
 AND2x2_ASAP7_75t_SL _220_ (.A(net73),
    .B(_033_),
    .Y(_112_));
 AO21x1_ASAP7_75t_SL _221_ (.A1(_078_),
    .A2(_032_),
    .B(_112_),
    .Y(_113_));
 AND3x1_ASAP7_75t_SL _222_ (.A(net76),
    .B(_000_),
    .C(_113_),
    .Y(_114_));
 AND2x2_ASAP7_75t_SL _223_ (.A(net73),
    .B(_029_),
    .Y(_115_));
 AO21x1_ASAP7_75t_SL _224_ (.A1(_078_),
    .A2(_028_),
    .B(_115_),
    .Y(_116_));
 AND2x2_ASAP7_75t_SL _225_ (.A(net74),
    .B(_027_),
    .Y(_117_));
 AO21x1_ASAP7_75t_SL _226_ (.A1(_078_),
    .A2(_026_),
    .B(_117_),
    .Y(_118_));
 AO22x1_ASAP7_75t_SL _227_ (.A1(_086_),
    .A2(_116_),
    .B1(_118_),
    .B2(_089_),
    .Y(_119_));
 AND2x2_ASAP7_75t_SL _228_ (.A(net80),
    .B(_031_),
    .Y(_120_));
 AO21x1_ASAP7_75t_SL _229_ (.A1(_078_),
    .A2(_030_),
    .B(_120_),
    .Y(_121_));
 AND3x1_ASAP7_75t_SL _230_ (.A(_093_),
    .B(_000_),
    .C(_121_),
    .Y(_122_));
 OR5x1_ASAP7_75t_SL _231_ (.A(_098_),
    .B(_111_),
    .C(_114_),
    .D(_119_),
    .E(_122_),
    .Y(_123_));
 AND2x2_ASAP7_75t_SL _232_ (.A(net80),
    .B(_025_),
    .Y(_124_));
 AO21x1_ASAP7_75t_SL _233_ (.A1(_078_),
    .A2(_024_),
    .B(_124_),
    .Y(_125_));
 AND3x1_ASAP7_75t_SL _234_ (.A(net76),
    .B(_000_),
    .C(_125_),
    .Y(_126_));
 AND2x2_ASAP7_75t_SL _235_ (.A(net74),
    .B(_021_),
    .Y(_127_));
 AO21x1_ASAP7_75t_SL _236_ (.A1(_078_),
    .A2(_020_),
    .B(_127_),
    .Y(_128_));
 AND2x2_ASAP7_75t_SL _237_ (.A(net74),
    .B(_019_),
    .Y(_129_));
 AO21x1_ASAP7_75t_SL _238_ (.A1(_078_),
    .A2(_018_),
    .B(_129_),
    .Y(_130_));
 AO22x1_ASAP7_75t_SL _239_ (.A1(_086_),
    .A2(_128_),
    .B1(_130_),
    .B2(_089_),
    .Y(_131_));
 AND2x2_ASAP7_75t_SL _240_ (.A(net80),
    .B(_023_),
    .Y(_132_));
 AO21x1_ASAP7_75t_SL _241_ (.A1(_078_),
    .A2(_022_),
    .B(_132_),
    .Y(_133_));
 AND3x1_ASAP7_75t_SL _242_ (.A(_093_),
    .B(_000_),
    .C(_133_),
    .Y(_134_));
 OR5x1_ASAP7_75t_SL _243_ (.A(_035_),
    .B(_111_),
    .C(_126_),
    .D(_131_),
    .E(_134_),
    .Y(_135_));
 AND4x1_ASAP7_75t_SL _244_ (.A(_097_),
    .B(_110_),
    .C(_123_),
    .D(_135_),
    .Y(_136_));
 NOR2x1_ASAP7_75t_SL _245_ (.A(_075_),
    .B(_136_),
    .Y(net35));
 BUFx4_ASAP7_75t_SL clkbuf_0_clock (.A(clock),
    .Y(clknet_0_clock));
 TAPCELL_ASAP7_75t_SL PHY_6 ();
 TAPCELL_ASAP7_75t_SL PHY_5 ();
 NOR2x1_ASAP7_75t_SL _249_ (.A(_033_),
    .B(net34),
    .Y(_139_));
 AO21x1_ASAP7_75t_SL _250_ (.A1(net1),
    .A2(net34),
    .B(_139_),
    .Y(_043_));
 TAPCELL_ASAP7_75t_SL PHY_4 ();
 NOR2x1_ASAP7_75t_SL _252_ (.A(_032_),
    .B(net34),
    .Y(_141_));
 AO21x1_ASAP7_75t_SL _253_ (.A1(net34),
    .A2(net12),
    .B(_141_),
    .Y(_044_));
 NOR2x1_ASAP7_75t_SL _254_ (.A(_031_),
    .B(net34),
    .Y(_142_));
 AO21x1_ASAP7_75t_SL _255_ (.A1(net34),
    .A2(net23),
    .B(_142_),
    .Y(_045_));
 NOR2x1_ASAP7_75t_SL _256_ (.A(_030_),
    .B(net34),
    .Y(_143_));
 AO21x1_ASAP7_75t_SL _257_ (.A1(net34),
    .A2(net26),
    .B(_143_),
    .Y(_046_));
 NOR2x1_ASAP7_75t_SL _258_ (.A(_029_),
    .B(net34),
    .Y(_144_));
 AO21x1_ASAP7_75t_SL _259_ (.A1(net34),
    .A2(net27),
    .B(_144_),
    .Y(_047_));
 NOR2x1_ASAP7_75t_SL _260_ (.A(_028_),
    .B(net34),
    .Y(_145_));
 AO21x1_ASAP7_75t_SL _261_ (.A1(net34),
    .A2(net28),
    .B(_145_),
    .Y(_048_));
 NOR2x1_ASAP7_75t_SL _262_ (.A(_027_),
    .B(net34),
    .Y(_146_));
 AO21x1_ASAP7_75t_SL _263_ (.A1(net34),
    .A2(net29),
    .B(_146_),
    .Y(_049_));
 NOR2x1_ASAP7_75t_SL _264_ (.A(_026_),
    .B(net34),
    .Y(_147_));
 AO21x1_ASAP7_75t_SL _265_ (.A1(net34),
    .A2(net30),
    .B(_147_),
    .Y(_050_));
 TAPCELL_ASAP7_75t_SL PHY_3 ();
 NOR2x1_ASAP7_75t_SL _267_ (.A(_025_),
    .B(net34),
    .Y(_149_));
 AO21x1_ASAP7_75t_SL _268_ (.A1(net34),
    .A2(net31),
    .B(_149_),
    .Y(_051_));
 NOR2x1_ASAP7_75t_SL _269_ (.A(_024_),
    .B(net34),
    .Y(_150_));
 AO21x1_ASAP7_75t_SL _270_ (.A1(net34),
    .A2(net32),
    .B(_150_),
    .Y(_052_));
 NOR2x1_ASAP7_75t_SL _271_ (.A(_023_),
    .B(net34),
    .Y(_151_));
 AO21x1_ASAP7_75t_SL _272_ (.A1(net34),
    .A2(net2),
    .B(_151_),
    .Y(_053_));
 TAPCELL_ASAP7_75t_SL PHY_2 ();
 NOR2x1_ASAP7_75t_SL _274_ (.A(_022_),
    .B(net34),
    .Y(_153_));
 AO21x1_ASAP7_75t_SL _275_ (.A1(net34),
    .A2(net3),
    .B(_153_),
    .Y(_054_));
 NOR2x1_ASAP7_75t_SL _276_ (.A(_021_),
    .B(net34),
    .Y(_154_));
 AO21x1_ASAP7_75t_SL _277_ (.A1(net34),
    .A2(net4),
    .B(_154_),
    .Y(_055_));
 NOR2x1_ASAP7_75t_SL _278_ (.A(_020_),
    .B(net34),
    .Y(_155_));
 AO21x1_ASAP7_75t_SL _279_ (.A1(net34),
    .A2(net5),
    .B(_155_),
    .Y(_056_));
 NOR2x1_ASAP7_75t_SL _280_ (.A(_019_),
    .B(net34),
    .Y(_156_));
 AO21x1_ASAP7_75t_SL _281_ (.A1(net34),
    .A2(net6),
    .B(_156_),
    .Y(_057_));
 NOR2x1_ASAP7_75t_SL _282_ (.A(_018_),
    .B(net34),
    .Y(_157_));
 AO21x1_ASAP7_75t_SL _283_ (.A1(net34),
    .A2(net7),
    .B(_157_),
    .Y(_058_));
 NOR2x1_ASAP7_75t_SL _284_ (.A(_017_),
    .B(net34),
    .Y(_158_));
 AO21x1_ASAP7_75t_SL _285_ (.A1(net34),
    .A2(net8),
    .B(_158_),
    .Y(_059_));
 NOR2x1_ASAP7_75t_SL _286_ (.A(_016_),
    .B(net34),
    .Y(_159_));
 AO21x1_ASAP7_75t_SL _287_ (.A1(net34),
    .A2(net9),
    .B(_159_),
    .Y(_060_));
 TAPCELL_ASAP7_75t_SL PHY_1 ();
 NOR2x1_ASAP7_75t_SL _289_ (.A(_015_),
    .B(net34),
    .Y(_161_));
 AO21x1_ASAP7_75t_SL _290_ (.A1(net34),
    .A2(net10),
    .B(_161_),
    .Y(_061_));
 NOR2x1_ASAP7_75t_SL _291_ (.A(_014_),
    .B(net34),
    .Y(_162_));
 AO21x1_ASAP7_75t_SL _292_ (.A1(net34),
    .A2(net11),
    .B(_162_),
    .Y(_062_));
 NOR2x1_ASAP7_75t_SL _293_ (.A(_013_),
    .B(net34),
    .Y(_163_));
 AO21x1_ASAP7_75t_SL _294_ (.A1(net34),
    .A2(net13),
    .B(_163_),
    .Y(_063_));
 TAPCELL_ASAP7_75t_SL PHY_0 ();
 NOR2x1_ASAP7_75t_SL _296_ (.A(_012_),
    .B(net34),
    .Y(_165_));
 AO21x1_ASAP7_75t_SL _297_ (.A1(net34),
    .A2(net14),
    .B(_165_),
    .Y(_064_));
 NOR2x1_ASAP7_75t_SL _298_ (.A(_011_),
    .B(net34),
    .Y(_166_));
 AO21x1_ASAP7_75t_SL _299_ (.A1(net34),
    .A2(net15),
    .B(_166_),
    .Y(_065_));
 NOR2x1_ASAP7_75t_SL _300_ (.A(_010_),
    .B(net34),
    .Y(_167_));
 AO21x1_ASAP7_75t_SL _301_ (.A1(net34),
    .A2(net16),
    .B(_167_),
    .Y(_066_));
 NOR2x1_ASAP7_75t_SL _302_ (.A(_009_),
    .B(net34),
    .Y(_168_));
 AO21x1_ASAP7_75t_SL _303_ (.A1(net34),
    .A2(net17),
    .B(_168_),
    .Y(_067_));
 NOR2x1_ASAP7_75t_SL _304_ (.A(_008_),
    .B(net34),
    .Y(_169_));
 AO21x1_ASAP7_75t_SL _305_ (.A1(net34),
    .A2(net18),
    .B(_169_),
    .Y(_068_));
 NOR2x1_ASAP7_75t_SL _306_ (.A(_007_),
    .B(net34),
    .Y(_170_));
 AO21x1_ASAP7_75t_SL _307_ (.A1(net34),
    .A2(net19),
    .B(_170_),
    .Y(_069_));
 NOR2x1_ASAP7_75t_SL _308_ (.A(_006_),
    .B(net34),
    .Y(_171_));
 AO21x1_ASAP7_75t_SL _309_ (.A1(net34),
    .A2(net20),
    .B(_171_),
    .Y(_070_));
 NOR2x1_ASAP7_75t_SL _310_ (.A(_005_),
    .B(net34),
    .Y(_172_));
 AO21x1_ASAP7_75t_SL _311_ (.A1(net34),
    .A2(net21),
    .B(_172_),
    .Y(_071_));
 NOR2x1_ASAP7_75t_SL _312_ (.A(_004_),
    .B(net34),
    .Y(_173_));
 AO21x1_ASAP7_75t_SL _313_ (.A1(net34),
    .A2(net22),
    .B(_173_),
    .Y(_072_));
 NOR2x1_ASAP7_75t_SL _314_ (.A(_003_),
    .B(net34),
    .Y(_174_));
 AO21x1_ASAP7_75t_SL _315_ (.A1(net34),
    .A2(net24),
    .B(_174_),
    .Y(_073_));
 NOR2x1_ASAP7_75t_SL _316_ (.A(_002_),
    .B(net34),
    .Y(_175_));
 AO21x1_ASAP7_75t_SL _317_ (.A1(net34),
    .A2(net25),
    .B(_175_),
    .Y(_074_));
 INVx2_ASAP7_75t_SL _318_ (.A(net34),
    .Y(_176_));
 AND2x2_ASAP7_75t_SL _319_ (.A(net74),
    .B(_176_),
    .Y(_038_));
 XOR2x1_ASAP7_75t_SL _320_ (.A(net75),
    .Y(_177_),
    .B(net77));
 AND2x2_ASAP7_75t_SL _321_ (.A(_176_),
    .B(_177_),
    .Y(_039_));
 OR3x1_ASAP7_75t_SL _322_ (.A(_001_),
    .B(_036_),
    .C(_000_),
    .Y(_178_));
 AO21x1_ASAP7_75t_SL _323_ (.A1(_078_),
    .A2(_093_),
    .B(_085_),
    .Y(_179_));
 AND3x1_ASAP7_75t_SL _324_ (.A(_176_),
    .B(_178_),
    .C(_179_),
    .Y(_040_));
 OR2x2_ASAP7_75t_SL _325_ (.A(_035_),
    .B(_178_),
    .Y(_180_));
 NAND2x1_ASAP7_75t_SL _326_ (.A(_035_),
    .B(net79),
    .Y(_181_));
 AND3x1_ASAP7_75t_SL _327_ (.A(_176_),
    .B(net81),
    .C(_181_),
    .Y(_041_));
 XNOR2x1_ASAP7_75t_SL _328_ (.B(_180_),
    .Y(_182_),
    .A(_111_));
 AND2x2_ASAP7_75t_SL _329_ (.A(_176_),
    .B(_182_),
    .Y(_042_));
 DFFLQNx1_ASAP7_75t_SL _330_ (.CLK(net72),
    .D(_038_),
    .QN(_001_));
 DFFLQNx1_ASAP7_75t_SL _331_ (.CLK(net71),
    .D(_039_),
    .QN(_036_));
 DFFLQNx1_ASAP7_75t_SL _332_ (.CLK(net70),
    .D(_040_),
    .QN(_000_));
 DFFLQNx1_ASAP7_75t_SL _333_ (.CLK(net69),
    .D(_041_),
    .QN(_035_));
 DFFLQNx1_ASAP7_75t_SL _334_ (.CLK(net68),
    .D(_042_),
    .QN(_034_));
 DFFLQNx1_ASAP7_75t_SL _335_ (.CLK(net67),
    .D(_043_),
    .QN(_033_));
 DFFLQNx1_ASAP7_75t_SL _336_ (.CLK(net66),
    .D(_044_),
    .QN(_032_));
 DFFLQNx1_ASAP7_75t_SL _337_ (.CLK(net65),
    .D(_045_),
    .QN(_031_));
 DFFLQNx1_ASAP7_75t_SL _338_ (.CLK(net64),
    .D(_046_),
    .QN(_030_));
 DFFLQNx1_ASAP7_75t_SL _339_ (.CLK(net63),
    .D(_047_),
    .QN(_029_));
 DFFLQNx1_ASAP7_75t_SL _340_ (.CLK(net62),
    .D(_048_),
    .QN(_028_));
 DFFLQNx1_ASAP7_75t_SL _341_ (.CLK(net61),
    .D(_049_),
    .QN(_027_));
 DFFLQNx1_ASAP7_75t_SL _342_ (.CLK(net60),
    .D(_050_),
    .QN(_026_));
 DFFLQNx1_ASAP7_75t_SL _343_ (.CLK(net59),
    .D(_051_),
    .QN(_025_));
 DFFLQNx1_ASAP7_75t_SL _344_ (.CLK(net58),
    .D(_052_),
    .QN(_024_));
 DFFLQNx1_ASAP7_75t_SL _345_ (.CLK(net57),
    .D(_053_),
    .QN(_023_));
 DFFLQNx1_ASAP7_75t_SL _346_ (.CLK(net56),
    .D(_054_),
    .QN(_022_));
 DFFLQNx1_ASAP7_75t_SL _347_ (.CLK(net55),
    .D(_055_),
    .QN(_021_));
 DFFLQNx1_ASAP7_75t_SL _348_ (.CLK(net54),
    .D(_056_),
    .QN(_020_));
 DFFLQNx1_ASAP7_75t_SL _349_ (.CLK(net53),
    .D(_057_),
    .QN(_019_));
 DFFLQNx1_ASAP7_75t_SL _350_ (.CLK(net52),
    .D(_058_),
    .QN(_018_));
 DFFLQNx1_ASAP7_75t_SL _351_ (.CLK(net51),
    .D(_059_),
    .QN(_017_));
 DFFLQNx1_ASAP7_75t_SL _352_ (.CLK(net50),
    .D(_060_),
    .QN(_016_));
 DFFLQNx1_ASAP7_75t_SL _353_ (.CLK(net49),
    .D(_061_),
    .QN(_015_));
 DFFLQNx1_ASAP7_75t_SL _354_ (.CLK(net48),
    .D(_062_),
    .QN(_014_));
 DFFLQNx1_ASAP7_75t_SL _355_ (.CLK(net47),
    .D(_063_),
    .QN(_013_));
 DFFLQNx1_ASAP7_75t_SL _356_ (.CLK(net46),
    .D(_064_),
    .QN(_012_));
 DFFLQNx1_ASAP7_75t_SL _357_ (.CLK(net45),
    .D(_065_),
    .QN(_011_));
 DFFLQNx1_ASAP7_75t_SL _358_ (.CLK(net44),
    .D(_066_),
    .QN(_010_));
 DFFLQNx1_ASAP7_75t_SL _359_ (.CLK(net43),
    .D(_067_),
    .QN(_009_));
 DFFLQNx1_ASAP7_75t_SL _360_ (.CLK(net42),
    .D(_068_),
    .QN(_008_));
 DFFLQNx1_ASAP7_75t_SL _361_ (.CLK(net41),
    .D(_069_),
    .QN(_007_));
 DFFLQNx1_ASAP7_75t_SL _362_ (.CLK(net40),
    .D(_070_),
    .QN(_006_));
 DFFLQNx1_ASAP7_75t_SL _363_ (.CLK(net39),
    .D(_071_),
    .QN(_005_));
 DFFLQNx1_ASAP7_75t_SL _364_ (.CLK(net38),
    .D(_072_),
    .QN(_004_));
 DFFLQNx1_ASAP7_75t_SL _365_ (.CLK(net37),
    .D(_073_),
    .QN(_003_));
 DFFLQNx1_ASAP7_75t_SL _366_ (.CLK(net36),
    .D(_074_),
    .QN(_002_));
 TAPCELL_ASAP7_75t_SL PHY_12 ();
 TAPCELL_ASAP7_75t_SL PHY_13 ();
 TAPCELL_ASAP7_75t_SL PHY_14 ();
 TAPCELL_ASAP7_75t_SL PHY_15 ();
 TAPCELL_ASAP7_75t_SL PHY_16 ();
 TAPCELL_ASAP7_75t_SL PHY_17 ();
 TAPCELL_ASAP7_75t_SL PHY_18 ();
 TAPCELL_ASAP7_75t_SL PHY_19 ();
 TAPCELL_ASAP7_75t_SL PHY_20 ();
 TAPCELL_ASAP7_75t_SL PHY_21 ();
 TAPCELL_ASAP7_75t_SL PHY_22 ();
 TAPCELL_ASAP7_75t_SL PHY_23 ();
 TAPCELL_ASAP7_75t_SL PHY_24 ();
 TAPCELL_ASAP7_75t_SL PHY_25 ();
 TAPCELL_ASAP7_75t_SL PHY_26 ();
 TAPCELL_ASAP7_75t_SL PHY_27 ();
 TAPCELL_ASAP7_75t_SL PHY_28 ();
 TAPCELL_ASAP7_75t_SL PHY_29 ();
 TAPCELL_ASAP7_75t_SL PHY_30 ();
 TAPCELL_ASAP7_75t_SL PHY_31 ();
 TAPCELL_ASAP7_75t_SL PHY_32 ();
 TAPCELL_ASAP7_75t_SL PHY_33 ();
 TAPCELL_ASAP7_75t_SL PHY_34 ();
 TAPCELL_ASAP7_75t_SL PHY_35 ();
 TAPCELL_ASAP7_75t_SL PHY_36 ();
 TAPCELL_ASAP7_75t_SL PHY_37 ();
 TAPCELL_ASAP7_75t_SL PHY_38 ();
 TAPCELL_ASAP7_75t_SL PHY_39 ();
 TAPCELL_ASAP7_75t_SL PHY_40 ();
 TAPCELL_ASAP7_75t_SL PHY_41 ();
 TAPCELL_ASAP7_75t_SL PHY_42 ();
 TAPCELL_ASAP7_75t_SL PHY_43 ();
 TAPCELL_ASAP7_75t_SL PHY_44 ();
 TAPCELL_ASAP7_75t_SL PHY_45 ();
 TAPCELL_ASAP7_75t_SL PHY_46 ();
 TAPCELL_ASAP7_75t_SL PHY_47 ();
 TAPCELL_ASAP7_75t_SL PHY_48 ();
 TAPCELL_ASAP7_75t_SL PHY_49 ();
 TAPCELL_ASAP7_75t_SL PHY_50 ();
 TAPCELL_ASAP7_75t_SL PHY_51 ();
 TAPCELL_ASAP7_75t_SL PHY_52 ();
 TAPCELL_ASAP7_75t_SL PHY_53 ();
 TAPCELL_ASAP7_75t_SL PHY_54 ();
 TAPCELL_ASAP7_75t_SL PHY_55 ();
 TAPCELL_ASAP7_75t_SL PHY_56 ();
 TAPCELL_ASAP7_75t_SL PHY_57 ();
 TAPCELL_ASAP7_75t_SL PHY_58 ();
 TAPCELL_ASAP7_75t_SL PHY_59 ();
 TAPCELL_ASAP7_75t_SL PHY_60 ();
 TAPCELL_ASAP7_75t_SL PHY_61 ();
 TAPCELL_ASAP7_75t_SL PHY_62 ();
 TAPCELL_ASAP7_75t_SL PHY_63 ();
 TAPCELL_ASAP7_75t_SL PHY_64 ();
 TAPCELL_ASAP7_75t_SL PHY_65 ();
 TAPCELL_ASAP7_75t_SL PHY_66 ();
 TAPCELL_ASAP7_75t_SL PHY_67 ();
 TAPCELL_ASAP7_75t_SL PHY_68 ();
 TAPCELL_ASAP7_75t_SL PHY_69 ();
 TAPCELL_ASAP7_75t_SL PHY_70 ();
 TAPCELL_ASAP7_75t_SL PHY_71 ();
 TAPCELL_ASAP7_75t_SL PHY_72 ();
 TAPCELL_ASAP7_75t_SL PHY_73 ();
 TAPCELL_ASAP7_75t_SL PHY_74 ();
 TAPCELL_ASAP7_75t_SL PHY_75 ();
 TAPCELL_ASAP7_75t_SL PHY_76 ();
 TAPCELL_ASAP7_75t_SL PHY_77 ();
 TAPCELL_ASAP7_75t_SL PHY_78 ();
 TAPCELL_ASAP7_75t_SL PHY_79 ();
 TAPCELL_ASAP7_75t_SL PHY_80 ();
 TAPCELL_ASAP7_75t_SL PHY_81 ();
 TAPCELL_ASAP7_75t_SL PHY_82 ();
 TAPCELL_ASAP7_75t_SL PHY_83 ();
 TAPCELL_ASAP7_75t_SL PHY_84 ();
 TAPCELL_ASAP7_75t_SL PHY_85 ();
 TAPCELL_ASAP7_75t_SL PHY_86 ();
 TAPCELL_ASAP7_75t_SL PHY_87 ();
 TAPCELL_ASAP7_75t_SL PHY_88 ();
 TAPCELL_ASAP7_75t_SL PHY_89 ();
 TAPCELL_ASAP7_75t_SL PHY_90 ();
 TAPCELL_ASAP7_75t_SL PHY_91 ();
 TAPCELL_ASAP7_75t_SL PHY_92 ();
 TAPCELL_ASAP7_75t_SL PHY_93 ();
 TAPCELL_ASAP7_75t_SL PHY_94 ();
 TAPCELL_ASAP7_75t_SL PHY_95 ();
 TAPCELL_ASAP7_75t_SL PHY_96 ();
 TAPCELL_ASAP7_75t_SL PHY_97 ();
 TAPCELL_ASAP7_75t_SL PHY_98 ();
 TAPCELL_ASAP7_75t_SL PHY_99 ();
 TAPCELL_ASAP7_75t_SL PHY_100 ();
 TAPCELL_ASAP7_75t_SL PHY_101 ();
 TAPCELL_ASAP7_75t_SL PHY_102 ();
 TAPCELL_ASAP7_75t_SL PHY_103 ();
 TAPCELL_ASAP7_75t_SL PHY_104 ();
 TAPCELL_ASAP7_75t_SL PHY_105 ();
 TAPCELL_ASAP7_75t_SL PHY_106 ();
 TAPCELL_ASAP7_75t_SL PHY_107 ();
 TAPCELL_ASAP7_75t_SL PHY_108 ();
 TAPCELL_ASAP7_75t_SL PHY_109 ();
 TAPCELL_ASAP7_75t_SL PHY_110 ();
 TAPCELL_ASAP7_75t_SL PHY_111 ();
 BUFx2_ASAP7_75t_SL input1 (.A(din[0]),
    .Y(net1));
 BUFx2_ASAP7_75t_SL input2 (.A(din[10]),
    .Y(net2));
 BUFx2_ASAP7_75t_SL input3 (.A(din[11]),
    .Y(net3));
 BUFx2_ASAP7_75t_SL input4 (.A(din[12]),
    .Y(net4));
 BUFx2_ASAP7_75t_SL input5 (.A(din[13]),
    .Y(net5));
 BUFx2_ASAP7_75t_SL input6 (.A(din[14]),
    .Y(net6));
 BUFx2_ASAP7_75t_SL input7 (.A(din[15]),
    .Y(net7));
 BUFx2_ASAP7_75t_SL input8 (.A(din[16]),
    .Y(net8));
 BUFx2_ASAP7_75t_SL input9 (.A(din[17]),
    .Y(net9));
 BUFx2_ASAP7_75t_SL input10 (.A(din[18]),
    .Y(net10));
 BUFx2_ASAP7_75t_SL input11 (.A(din[19]),
    .Y(net11));
 BUFx2_ASAP7_75t_SL input12 (.A(din[1]),
    .Y(net12));
 BUFx2_ASAP7_75t_SL input13 (.A(din[20]),
    .Y(net13));
 BUFx2_ASAP7_75t_SL input14 (.A(din[21]),
    .Y(net14));
 BUFx2_ASAP7_75t_SL input15 (.A(din[22]),
    .Y(net15));
 BUFx2_ASAP7_75t_SL input16 (.A(din[23]),
    .Y(net16));
 BUFx2_ASAP7_75t_SL input17 (.A(din[24]),
    .Y(net17));
 BUFx2_ASAP7_75t_SL input18 (.A(din[25]),
    .Y(net18));
 BUFx2_ASAP7_75t_SL input19 (.A(din[26]),
    .Y(net19));
 BUFx2_ASAP7_75t_SL input20 (.A(din[27]),
    .Y(net20));
 BUFx2_ASAP7_75t_SL input21 (.A(din[28]),
    .Y(net21));
 BUFx2_ASAP7_75t_SL input22 (.A(din[29]),
    .Y(net22));
 BUFx2_ASAP7_75t_SL input23 (.A(din[2]),
    .Y(net23));
 BUFx2_ASAP7_75t_SL input24 (.A(din[30]),
    .Y(net24));
 BUFx2_ASAP7_75t_SL input25 (.A(din[31]),
    .Y(net25));
 BUFx2_ASAP7_75t_SL input26 (.A(din[3]),
    .Y(net26));
 BUFx2_ASAP7_75t_SL input27 (.A(din[4]),
    .Y(net27));
 BUFx2_ASAP7_75t_SL input28 (.A(din[5]),
    .Y(net28));
 BUFx2_ASAP7_75t_SL input29 (.A(din[6]),
    .Y(net29));
 BUFx2_ASAP7_75t_SL input30 (.A(din[7]),
    .Y(net30));
 BUFx2_ASAP7_75t_SL input31 (.A(din[8]),
    .Y(net31));
 BUFx2_ASAP7_75t_SL input32 (.A(din[9]),
    .Y(net32));
 BUFx2_ASAP7_75t_SL input33 (.A(enable),
    .Y(net33));
 BUFx16f_ASAP7_75t_SL input34 (.A(load),
    .Y(net34));
 BUFx2_ASAP7_75t_SL output35 (.A(net35),
    .Y(dout));
 INVx1_ASAP7_75t_SL _246__1 (.A(clknet_2_1__leaf_clock),
    .Y(net36));
 INVx1_ASAP7_75t_SL _246__2 (.A(clknet_2_1__leaf_clock),
    .Y(net37));
 INVx1_ASAP7_75t_SL _246__3 (.A(clknet_2_1__leaf_clock),
    .Y(net38));
 INVx1_ASAP7_75t_SL _246__4 (.A(clknet_2_1__leaf_clock),
    .Y(net39));
 INVx1_ASAP7_75t_SL _246__5 (.A(clknet_2_3__leaf_clock),
    .Y(net40));
 INVx1_ASAP7_75t_SL _246__6 (.A(clknet_2_3__leaf_clock),
    .Y(net41));
 INVx1_ASAP7_75t_SL _246__7 (.A(clknet_2_2__leaf_clock),
    .Y(net42));
 INVx1_ASAP7_75t_SL _246__8 (.A(clknet_2_2__leaf_clock),
    .Y(net43));
 INVx1_ASAP7_75t_SL _246__9 (.A(clknet_2_2__leaf_clock),
    .Y(net44));
 INVx1_ASAP7_75t_SL _246__10 (.A(clknet_2_2__leaf_clock),
    .Y(net45));
 INVx1_ASAP7_75t_SL _246__11 (.A(clknet_2_0__leaf_clock),
    .Y(net46));
 INVx1_ASAP7_75t_SL _246__12 (.A(clknet_2_0__leaf_clock),
    .Y(net47));
 INVx1_ASAP7_75t_SL _246__13 (.A(clknet_2_2__leaf_clock),
    .Y(net48));
 INVx1_ASAP7_75t_SL _246__14 (.A(clknet_2_2__leaf_clock),
    .Y(net49));
 INVx1_ASAP7_75t_SL _246__15 (.A(clknet_2_2__leaf_clock),
    .Y(net50));
 INVx1_ASAP7_75t_SL _246__16 (.A(clknet_2_2__leaf_clock),
    .Y(net51));
 INVx1_ASAP7_75t_SL _246__17 (.A(clknet_2_0__leaf_clock),
    .Y(net52));
 INVx1_ASAP7_75t_SL _246__18 (.A(clknet_2_0__leaf_clock),
    .Y(net53));
 INVx1_ASAP7_75t_SL _246__19 (.A(clknet_2_0__leaf_clock),
    .Y(net54));
 INVx1_ASAP7_75t_SL _246__20 (.A(clknet_2_0__leaf_clock),
    .Y(net55));
 INVx1_ASAP7_75t_SL _246__21 (.A(clknet_2_3__leaf_clock),
    .Y(net56));
 INVx1_ASAP7_75t_SL _246__22 (.A(clknet_2_3__leaf_clock),
    .Y(net57));
 INVx1_ASAP7_75t_SL _246__23 (.A(clknet_2_3__leaf_clock),
    .Y(net58));
 INVx1_ASAP7_75t_SL _246__24 (.A(clknet_2_1__leaf_clock),
    .Y(net59));
 INVx1_ASAP7_75t_SL _246__25 (.A(clknet_2_1__leaf_clock),
    .Y(net60));
 INVx1_ASAP7_75t_SL _246__26 (.A(clknet_2_1__leaf_clock),
    .Y(net61));
 INVx1_ASAP7_75t_SL _246__27 (.A(clknet_2_0__leaf_clock),
    .Y(net62));
 INVx1_ASAP7_75t_SL _246__28 (.A(clknet_2_0__leaf_clock),
    .Y(net63));
 INVx1_ASAP7_75t_SL _246__29 (.A(clknet_2_3__leaf_clock),
    .Y(net64));
 INVx1_ASAP7_75t_SL _246__30 (.A(clknet_2_3__leaf_clock),
    .Y(net65));
 INVx1_ASAP7_75t_SL _246__31 (.A(clknet_2_3__leaf_clock),
    .Y(net66));
 INVx1_ASAP7_75t_SL _246__32 (.A(clknet_2_3__leaf_clock),
    .Y(net67));
 INVx1_ASAP7_75t_SL _33 (.A(clknet_2_2__leaf_clock),
    .Y(net68));
 INVx1_ASAP7_75t_SL _33_34 (.A(clknet_2_2__leaf_clock),
    .Y(net69));
 INVx1_ASAP7_75t_SL _33_35 (.A(clknet_2_3__leaf_clock),
    .Y(net70));
 INVx1_ASAP7_75t_SL _33_36 (.A(clknet_2_1__leaf_clock),
    .Y(net71));
 INVx1_ASAP7_75t_SL _33_37 (.A(clknet_2_0__leaf_clock),
    .Y(net72));
 BUFx4_ASAP7_75t_SL clkbuf_2_0__f_clock (.A(clknet_0_clock),
    .Y(clknet_2_0__leaf_clock));
 BUFx4_ASAP7_75t_SL clkbuf_2_1__f_clock (.A(clknet_0_clock),
    .Y(clknet_2_1__leaf_clock));
 BUFx4_ASAP7_75t_SL clkbuf_2_2__f_clock (.A(clknet_0_clock),
    .Y(clknet_2_2__leaf_clock));
 BUFx4_ASAP7_75t_SL clkbuf_2_3__f_clock (.A(clknet_0_clock),
    .Y(clknet_2_3__leaf_clock));
 BUFx3_ASAP7_75t_SL split38 (.A(_001_),
    .Y(net73));
 BUFx4f_ASAP7_75t_SL rebuffer39 (.A(_001_),
    .Y(net74));
 BUFx2_ASAP7_75t_SL rebuffer40 (.A(net80),
    .Y(net75));
 BUFx2_ASAP7_75t_SL rebuffer41 (.A(_036_),
    .Y(net76));
 BUFx2_ASAP7_75t_SL rebuffer42 (.A(_036_),
    .Y(net77));
 BUFx2_ASAP7_75t_SL split43 (.A(_000_),
    .Y(net78));
 BUFx2_ASAP7_75t_SL rebuffer44 (.A(_178_),
    .Y(net79));
 BUFx2_ASAP7_75t_SL rebuffer45 (.A(_001_),
    .Y(net80));
 BUFx2_ASAP7_75t_SL rebuffer46 (.A(_180_),
    .Y(net81));
 DECAPx10_ASAP7_75t_SL FILLER_0_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_68 ();
 DECAPx6_ASAP7_75t_SL FILLER_0_90 ();
 DECAPx1_ASAP7_75t_SL FILLER_0_104 ();
 FILLERxp5_ASAP7_75t_SL FILLER_0_108 ();
 DECAPx6_ASAP7_75t_SL FILLER_0_114 ();
 FILLER_ASAP7_75t_SL FILLER_0_128 ();
 FILLER_ASAP7_75t_SL FILLER_0_135 ();
 DECAPx4_ASAP7_75t_SL FILLER_0_142 ();
 FILLER_ASAP7_75t_SL FILLER_0_152 ();
 DECAPx2_ASAP7_75t_SL FILLER_0_159 ();
 FILLER_ASAP7_75t_SL FILLER_0_165 ();
 DECAPx6_ASAP7_75t_SL FILLER_0_172 ();
 FILLERxp5_ASAP7_75t_SL FILLER_0_186 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_192 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_214 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_236 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_258 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_0_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_68 ();
 DECAPx6_ASAP7_75t_SL FILLER_1_90 ();
 DECAPx1_ASAP7_75t_SL FILLER_1_104 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_113 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_135 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_157 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_179 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_201 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_223 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_245 ();
 DECAPx6_ASAP7_75t_SL FILLER_1_267 ();
 FILLER_ASAP7_75t_SL FILLER_1_281 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_2_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_2_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_3_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_3_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_4_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_4_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_5_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_5_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_6_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_6_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_7_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_7_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_8_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_8_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_9_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_9_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_10_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_10_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_11_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_11_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_12_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_12_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_13_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_13_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_13_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_14_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_14_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_15_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_15_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_15_280 ();
 FILLER_ASAP7_75t_SL FILLER_16_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_9 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_31 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_53 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_75 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_97 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_119 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_141 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_163 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_185 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_207 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_229 ();
 DECAPx10_ASAP7_75t_SL FILLER_16_251 ();
 DECAPx4_ASAP7_75t_SL FILLER_16_273 ();
 DECAPx2_ASAP7_75t_SL FILLER_17_2 ();
 FILLER_ASAP7_75t_SL FILLER_17_8 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_16 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_38 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_60 ();
 DECAPx6_ASAP7_75t_SL FILLER_17_82 ();
 DECAPx1_ASAP7_75t_SL FILLER_17_96 ();
 DECAPx6_ASAP7_75t_SL FILLER_17_106 ();
 DECAPx2_ASAP7_75t_SL FILLER_17_120 ();
 FILLERxp5_ASAP7_75t_SL FILLER_17_126 ();
 FILLER_ASAP7_75t_SL FILLER_17_133 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_141 ();
 DECAPx6_ASAP7_75t_SL FILLER_17_163 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_17_177 ();
 FILLER_ASAP7_75t_SL FILLER_17_186 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_194 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_216 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_238 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_260 ();
 FILLERxp5_ASAP7_75t_SL FILLER_17_282 ();
 FILLER_ASAP7_75t_SL FILLER_18_2 ();
 FILLER_ASAP7_75t_SL FILLER_18_7 ();
 DECAPx1_ASAP7_75t_SL FILLER_18_29 ();
 FILLERxp5_ASAP7_75t_SL FILLER_18_33 ();
 DECAPx10_ASAP7_75t_SL FILLER_18_40 ();
 DECAPx10_ASAP7_75t_SL FILLER_18_62 ();
 DECAPx6_ASAP7_75t_SL FILLER_18_84 ();
 DECAPx1_ASAP7_75t_SL FILLER_18_98 ();
 FILLER_ASAP7_75t_SL FILLER_18_108 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_18_116 ();
 DECAPx1_ASAP7_75t_SL FILLER_18_139 ();
 DECAPx2_ASAP7_75t_SL FILLER_18_149 ();
 DECAPx2_ASAP7_75t_SL FILLER_18_161 ();
 DECAPx1_ASAP7_75t_SL FILLER_18_173 ();
 FILLERxp5_ASAP7_75t_SL FILLER_18_177 ();
 DECAPx10_ASAP7_75t_SL FILLER_18_198 ();
 DECAPx10_ASAP7_75t_SL FILLER_18_220 ();
 DECAPx2_ASAP7_75t_SL FILLER_18_242 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_18_248 ();
 DECAPx10_ASAP7_75t_SL FILLER_18_256 ();
 DECAPx1_ASAP7_75t_SL FILLER_18_278 ();
 FILLERxp5_ASAP7_75t_SL FILLER_18_282 ();
 FILLER_ASAP7_75t_SL FILLER_19_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_19_9 ();
 DECAPx10_ASAP7_75t_SL FILLER_19_32 ();
 DECAPx10_ASAP7_75t_SL FILLER_19_54 ();
 DECAPx6_ASAP7_75t_SL FILLER_19_76 ();
 DECAPx2_ASAP7_75t_SL FILLER_19_90 ();
 DECAPx1_ASAP7_75t_SL FILLER_19_116 ();
 FILLER_ASAP7_75t_SL FILLER_19_123 ();
 DECAPx2_ASAP7_75t_SL FILLER_19_145 ();
 FILLER_ASAP7_75t_SL FILLER_19_171 ();
 FILLER_ASAP7_75t_SL FILLER_19_179 ();
 FILLER_ASAP7_75t_SL FILLER_19_184 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_19_192 ();
 FILLER_ASAP7_75t_SL FILLER_19_201 ();
 DECAPx10_ASAP7_75t_SL FILLER_19_209 ();
 DECAPx10_ASAP7_75t_SL FILLER_19_231 ();
 DECAPx10_ASAP7_75t_SL FILLER_19_253 ();
 DECAPx2_ASAP7_75t_SL FILLER_19_275 ();
 FILLER_ASAP7_75t_SL FILLER_19_281 ();
 FILLER_ASAP7_75t_SL FILLER_20_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_20_9 ();
 DECAPx1_ASAP7_75t_SL FILLER_20_18 ();
 FILLERxp5_ASAP7_75t_SL FILLER_20_22 ();
 FILLER_ASAP7_75t_SL FILLER_20_29 ();
 FILLER_ASAP7_75t_SL FILLER_20_34 ();
 DECAPx10_ASAP7_75t_SL FILLER_20_42 ();
 DECAPx10_ASAP7_75t_SL FILLER_20_64 ();
 DECAPx4_ASAP7_75t_SL FILLER_20_86 ();
 FILLERxp5_ASAP7_75t_SL FILLER_20_96 ();
 FILLER_ASAP7_75t_SL FILLER_20_100 ();
 FILLER_ASAP7_75t_SL FILLER_20_122 ();
 DECAPx1_ASAP7_75t_SL FILLER_20_130 ();
 FILLERxp5_ASAP7_75t_SL FILLER_20_134 ();
 FILLER_ASAP7_75t_SL FILLER_20_141 ();
 DECAPx1_ASAP7_75t_SL FILLER_20_149 ();
 FILLER_ASAP7_75t_SL FILLER_20_173 ();
 DECAPx1_ASAP7_75t_SL FILLER_20_181 ();
 DECAPx10_ASAP7_75t_SL FILLER_20_205 ();
 DECAPx10_ASAP7_75t_SL FILLER_20_227 ();
 DECAPx10_ASAP7_75t_SL FILLER_20_249 ();
 DECAPx4_ASAP7_75t_SL FILLER_20_271 ();
 FILLER_ASAP7_75t_SL FILLER_20_281 ();
 DECAPx2_ASAP7_75t_SL FILLER_21_2 ();
 FILLER_ASAP7_75t_SL FILLER_21_8 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_21_16 ();
 DECAPx6_ASAP7_75t_SL FILLER_21_25 ();
 FILLER_ASAP7_75t_SL FILLER_21_39 ();
 DECAPx10_ASAP7_75t_SL FILLER_21_47 ();
 DECAPx10_ASAP7_75t_SL FILLER_21_69 ();
 DECAPx4_ASAP7_75t_SL FILLER_21_91 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_21_101 ();
 DECAPx2_ASAP7_75t_SL FILLER_21_107 ();
 FILLER_ASAP7_75t_SL FILLER_21_119 ();
 DECAPx2_ASAP7_75t_SL FILLER_21_127 ();
 DECAPx6_ASAP7_75t_SL FILLER_21_139 ();
 FILLER_ASAP7_75t_SL FILLER_21_153 ();
 FILLER_ASAP7_75t_SL FILLER_21_158 ();
 DECAPx2_ASAP7_75t_SL FILLER_21_163 ();
 FILLER_ASAP7_75t_SL FILLER_21_169 ();
 DECAPx2_ASAP7_75t_SL FILLER_21_177 ();
 FILLER_ASAP7_75t_SL FILLER_21_183 ();
 DECAPx4_ASAP7_75t_SL FILLER_21_191 ();
 FILLER_ASAP7_75t_SL FILLER_21_201 ();
 DECAPx10_ASAP7_75t_SL FILLER_21_206 ();
 DECAPx10_ASAP7_75t_SL FILLER_21_228 ();
 DECAPx10_ASAP7_75t_SL FILLER_21_250 ();
 DECAPx4_ASAP7_75t_SL FILLER_21_272 ();
 FILLERxp5_ASAP7_75t_SL FILLER_21_282 ();
 DECAPx2_ASAP7_75t_SL FILLER_22_2 ();
 FILLERxp5_ASAP7_75t_SL FILLER_22_8 ();
 DECAPx4_ASAP7_75t_SL FILLER_22_29 ();
 FILLER_ASAP7_75t_SL FILLER_22_45 ();
 DECAPx10_ASAP7_75t_SL FILLER_22_53 ();
 DECAPx10_ASAP7_75t_SL FILLER_22_75 ();
 DECAPx10_ASAP7_75t_SL FILLER_22_97 ();
 DECAPx2_ASAP7_75t_SL FILLER_22_119 ();
 FILLER_ASAP7_75t_SL FILLER_22_125 ();
 DECAPx10_ASAP7_75t_SL FILLER_22_130 ();
 DECAPx6_ASAP7_75t_SL FILLER_22_152 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_22_166 ();
 DECAPx4_ASAP7_75t_SL FILLER_22_175 ();
 FILLER_ASAP7_75t_SL FILLER_22_185 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_22_207 ();
 DECAPx10_ASAP7_75t_SL FILLER_22_216 ();
 DECAPx4_ASAP7_75t_SL FILLER_22_238 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_22_248 ();
 DECAPx10_ASAP7_75t_SL FILLER_22_256 ();
 DECAPx1_ASAP7_75t_SL FILLER_22_278 ();
 FILLERxp5_ASAP7_75t_SL FILLER_22_282 ();
 DECAPx2_ASAP7_75t_SL FILLER_23_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_23_8 ();
 DECAPx2_ASAP7_75t_SL FILLER_23_14 ();
 FILLER_ASAP7_75t_SL FILLER_23_20 ();
 DECAPx2_ASAP7_75t_SL FILLER_23_27 ();
 DECAPx10_ASAP7_75t_SL FILLER_23_53 ();
 DECAPx1_ASAP7_75t_SL FILLER_23_75 ();
 FILLERxp5_ASAP7_75t_SL FILLER_23_79 ();
 DECAPx10_ASAP7_75t_SL FILLER_23_104 ();
 DECAPx10_ASAP7_75t_SL FILLER_23_126 ();
 DECAPx10_ASAP7_75t_SL FILLER_23_148 ();
 DECAPx6_ASAP7_75t_SL FILLER_23_170 ();
 DECAPx1_ASAP7_75t_SL FILLER_23_184 ();
 FILLERxp5_ASAP7_75t_SL FILLER_23_188 ();
 DECAPx6_ASAP7_75t_SL FILLER_23_192 ();
 FILLERxp5_ASAP7_75t_SL FILLER_23_206 ();
 DECAPx10_ASAP7_75t_SL FILLER_23_213 ();
 DECAPx6_ASAP7_75t_SL FILLER_23_235 ();
 FILLER_ASAP7_75t_SL FILLER_23_249 ();
 DECAPx10_ASAP7_75t_SL FILLER_23_256 ();
 DECAPx1_ASAP7_75t_SL FILLER_23_278 ();
 FILLERxp5_ASAP7_75t_SL FILLER_23_282 ();
 FILLER_ASAP7_75t_SL FILLER_24_2 ();
 DECAPx1_ASAP7_75t_SL FILLER_24_9 ();
 FILLERxp5_ASAP7_75t_SL FILLER_24_13 ();
 FILLER_ASAP7_75t_SL FILLER_24_34 ();
 FILLER_ASAP7_75t_SL FILLER_24_42 ();
 DECAPx1_ASAP7_75t_SL FILLER_24_50 ();
 DECAPx10_ASAP7_75t_SL FILLER_24_63 ();
 DECAPx10_ASAP7_75t_SL FILLER_24_85 ();
 DECAPx6_ASAP7_75t_SL FILLER_24_107 ();
 DECAPx1_ASAP7_75t_SL FILLER_24_121 ();
 DECAPx1_ASAP7_75t_SL FILLER_24_134 ();
 FILLERxp5_ASAP7_75t_SL FILLER_24_138 ();
 DECAPx10_ASAP7_75t_SL FILLER_24_159 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_24_181 ();
 FILLER_ASAP7_75t_SL FILLER_24_204 ();
 DECAPx10_ASAP7_75t_SL FILLER_24_212 ();
 DECAPx10_ASAP7_75t_SL FILLER_24_234 ();
 DECAPx10_ASAP7_75t_SL FILLER_24_256 ();
 DECAPx1_ASAP7_75t_SL FILLER_24_278 ();
 FILLERxp5_ASAP7_75t_SL FILLER_24_282 ();
 DECAPx4_ASAP7_75t_SL FILLER_25_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_25_12 ();
 FILLER_ASAP7_75t_SL FILLER_25_21 ();
 DECAPx1_ASAP7_75t_SL FILLER_25_26 ();
 FILLERxp5_ASAP7_75t_SL FILLER_25_30 ();
 FILLER_ASAP7_75t_SL FILLER_25_37 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_45 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_67 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_89 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_25_111 ();
 FILLER_ASAP7_75t_SL FILLER_25_118 ();
 FILLER_ASAP7_75t_SL FILLER_25_140 ();
 FILLER_ASAP7_75t_SL FILLER_25_148 ();
 FILLER_ASAP7_75t_SL FILLER_25_153 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_158 ();
 DECAPx2_ASAP7_75t_SL FILLER_25_180 ();
 FILLER_ASAP7_75t_SL FILLER_25_192 ();
 FILLER_ASAP7_75t_SL FILLER_25_200 ();
 FILLER_ASAP7_75t_SL FILLER_25_208 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_213 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_235 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_257 ();
 DECAPx1_ASAP7_75t_SL FILLER_25_279 ();
 DECAPx2_ASAP7_75t_SL FILLER_26_2 ();
 FILLER_ASAP7_75t_SL FILLER_26_8 ();
 DECAPx1_ASAP7_75t_SL FILLER_26_30 ();
 FILLERxp5_ASAP7_75t_SL FILLER_26_34 ();
 DECAPx6_ASAP7_75t_SL FILLER_26_38 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_26_52 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_62 ();
 DECAPx6_ASAP7_75t_SL FILLER_26_84 ();
 FILLER_ASAP7_75t_SL FILLER_26_98 ();
 FILLER_ASAP7_75t_SL FILLER_26_106 ();
 FILLER_ASAP7_75t_SL FILLER_26_114 ();
 FILLER_ASAP7_75t_SL FILLER_26_122 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_26_130 ();
 FILLER_ASAP7_75t_SL FILLER_26_139 ();
 FILLER_ASAP7_75t_SL FILLER_26_153 ();
 FILLER_ASAP7_75t_SL FILLER_26_162 ();
 FILLER_ASAP7_75t_SL FILLER_26_170 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_26_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_26_280 ();
 FILLER_ASAP7_75t_SL FILLER_27_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_27_9 ();
 FILLER_ASAP7_75t_SL FILLER_27_15 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_27_23 ();
 DECAPx2_ASAP7_75t_SL FILLER_27_32 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_27_38 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_47 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_69 ();
 DECAPx1_ASAP7_75t_SL FILLER_27_91 ();
 FILLERxp5_ASAP7_75t_SL FILLER_27_95 ();
 FILLER_ASAP7_75t_SL FILLER_27_116 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_27_121 ();
 FILLER_ASAP7_75t_SL FILLER_27_130 ();
 FILLER_ASAP7_75t_SL FILLER_27_138 ();
 FILLER_ASAP7_75t_SL FILLER_27_145 ();
 FILLER_ASAP7_75t_SL FILLER_27_152 ();
 FILLER_ASAP7_75t_SL FILLER_27_157 ();
 FILLER_ASAP7_75t_SL FILLER_27_167 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_175 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_197 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_219 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_241 ();
 DECAPx6_ASAP7_75t_SL FILLER_27_263 ();
 DECAPx2_ASAP7_75t_SL FILLER_27_277 ();
 DECAPx2_ASAP7_75t_SL FILLER_28_2 ();
 FILLER_ASAP7_75t_SL FILLER_28_8 ();
 FILLER_ASAP7_75t_SL FILLER_28_16 ();
 DECAPx4_ASAP7_75t_SL FILLER_28_24 ();
 DECAPx2_ASAP7_75t_SL FILLER_28_40 ();
 FILLERxp5_ASAP7_75t_SL FILLER_28_46 ();
 FILLER_ASAP7_75t_SL FILLER_28_53 ();
 DECAPx10_ASAP7_75t_SL FILLER_28_64 ();
 DECAPx4_ASAP7_75t_SL FILLER_28_86 ();
 FILLER_ASAP7_75t_SL FILLER_28_96 ();
 DECAPx1_ASAP7_75t_SL FILLER_28_101 ();
 FILLER_ASAP7_75t_SL FILLER_28_117 ();
 DECAPx1_ASAP7_75t_SL FILLER_28_127 ();
 FILLERxp5_ASAP7_75t_SL FILLER_28_131 ();
 FILLER_ASAP7_75t_SL FILLER_28_138 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_28_144 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_28_155 ();
 FILLER_ASAP7_75t_SL FILLER_28_166 ();
 DECAPx6_ASAP7_75t_SL FILLER_28_175 ();
 FILLERxp5_ASAP7_75t_SL FILLER_28_189 ();
 DECAPx4_ASAP7_75t_SL FILLER_28_196 ();
 FILLERxp5_ASAP7_75t_SL FILLER_28_206 ();
 DECAPx10_ASAP7_75t_SL FILLER_28_213 ();
 DECAPx10_ASAP7_75t_SL FILLER_28_235 ();
 DECAPx10_ASAP7_75t_SL FILLER_28_257 ();
 DECAPx1_ASAP7_75t_SL FILLER_28_279 ();
 DECAPx2_ASAP7_75t_SL FILLER_29_2 ();
 FILLER_ASAP7_75t_SL FILLER_29_28 ();
 FILLER_ASAP7_75t_SL FILLER_29_50 ();
 FILLER_ASAP7_75t_SL FILLER_29_61 ();
 DECAPx10_ASAP7_75t_SL FILLER_29_70 ();
 DECAPx4_ASAP7_75t_SL FILLER_29_92 ();
 FILLER_ASAP7_75t_SL FILLER_29_122 ();
 FILLER_ASAP7_75t_SL FILLER_29_130 ();
 FILLER_ASAP7_75t_SL FILLER_29_138 ();
 FILLER_ASAP7_75t_SL FILLER_29_146 ();
 DECAPx1_ASAP7_75t_SL FILLER_29_155 ();
 FILLERxp5_ASAP7_75t_SL FILLER_29_159 ();
 FILLER_ASAP7_75t_SL FILLER_29_168 ();
 FILLER_ASAP7_75t_SL FILLER_29_176 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_29_184 ();
 FILLER_ASAP7_75t_SL FILLER_29_207 ();
 DECAPx10_ASAP7_75t_SL FILLER_29_215 ();
 DECAPx10_ASAP7_75t_SL FILLER_29_237 ();
 DECAPx1_ASAP7_75t_SL FILLER_29_259 ();
 FILLER_ASAP7_75t_SL FILLER_29_269 ();
 FILLER_ASAP7_75t_SL FILLER_29_274 ();
 FILLER_ASAP7_75t_SL FILLER_29_281 ();
 FILLER_ASAP7_75t_SL FILLER_30_2 ();
 FILLER_ASAP7_75t_SL FILLER_30_9 ();
 FILLER_ASAP7_75t_SL FILLER_30_16 ();
 DECAPx1_ASAP7_75t_SL FILLER_30_21 ();
 FILLER_ASAP7_75t_SL FILLER_30_30 ();
 DECAPx1_ASAP7_75t_SL FILLER_30_38 ();
 FILLERxp5_ASAP7_75t_SL FILLER_30_42 ();
 DECAPx10_ASAP7_75t_SL FILLER_30_49 ();
 DECAPx10_ASAP7_75t_SL FILLER_30_71 ();
 DECAPx4_ASAP7_75t_SL FILLER_30_93 ();
 FILLER_ASAP7_75t_SL FILLER_30_106 ();
 FILLER_ASAP7_75t_SL FILLER_30_115 ();
 FILLER_ASAP7_75t_SL FILLER_30_123 ();
 FILLER_ASAP7_75t_SL FILLER_30_130 ();
 DECAPx2_ASAP7_75t_SL FILLER_30_152 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_30_158 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_30_167 ();
 DECAPx10_ASAP7_75t_SL FILLER_30_176 ();
 DECAPx2_ASAP7_75t_SL FILLER_30_198 ();
 FILLERxp5_ASAP7_75t_SL FILLER_30_204 ();
 DECAPx10_ASAP7_75t_SL FILLER_30_208 ();
 DECAPx10_ASAP7_75t_SL FILLER_30_230 ();
 FILLERxp5_ASAP7_75t_SL FILLER_30_252 ();
 DECAPx2_ASAP7_75t_SL FILLER_30_258 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_30_264 ();
 DECAPx1_ASAP7_75t_SL FILLER_30_272 ();
 FILLER_ASAP7_75t_SL FILLER_30_281 ();
 DECAPx1_ASAP7_75t_SL FILLER_31_2 ();
 FILLERxp5_ASAP7_75t_SL FILLER_31_6 ();
 DECAPx1_ASAP7_75t_SL FILLER_31_27 ();
 FILLERxp5_ASAP7_75t_SL FILLER_31_31 ();
 DECAPx2_ASAP7_75t_SL FILLER_31_35 ();
 DECAPx10_ASAP7_75t_SL FILLER_31_47 ();
 DECAPx10_ASAP7_75t_SL FILLER_31_69 ();
 DECAPx6_ASAP7_75t_SL FILLER_31_91 ();
 FILLER_ASAP7_75t_SL FILLER_31_105 ();
 FILLER_ASAP7_75t_SL FILLER_31_113 ();
 FILLER_ASAP7_75t_SL FILLER_31_120 ();
 FILLER_ASAP7_75t_SL FILLER_31_127 ();
 FILLER_ASAP7_75t_SL FILLER_31_132 ();
 DECAPx6_ASAP7_75t_SL FILLER_31_137 ();
 FILLERxp5_ASAP7_75t_SL FILLER_31_151 ();
 DECAPx6_ASAP7_75t_SL FILLER_31_157 ();
 DECAPx1_ASAP7_75t_SL FILLER_31_171 ();
 FILLER_ASAP7_75t_SL FILLER_31_195 ();
 FILLER_ASAP7_75t_SL FILLER_31_203 ();
 DECAPx10_ASAP7_75t_SL FILLER_31_211 ();
 DECAPx10_ASAP7_75t_SL FILLER_31_233 ();
 DECAPx10_ASAP7_75t_SL FILLER_31_255 ();
 DECAPx2_ASAP7_75t_SL FILLER_31_277 ();
 DECAPx2_ASAP7_75t_SL FILLER_32_2 ();
 FILLER_ASAP7_75t_SL FILLER_32_14 ();
 FILLER_ASAP7_75t_SL FILLER_32_36 ();
 DECAPx10_ASAP7_75t_SL FILLER_32_44 ();
 DECAPx10_ASAP7_75t_SL FILLER_32_66 ();
 DECAPx10_ASAP7_75t_SL FILLER_32_88 ();
 DECAPx2_ASAP7_75t_SL FILLER_32_110 ();
 FILLERxp5_ASAP7_75t_SL FILLER_32_116 ();
 DECAPx10_ASAP7_75t_SL FILLER_32_122 ();
 DECAPx10_ASAP7_75t_SL FILLER_32_144 ();
 DECAPx10_ASAP7_75t_SL FILLER_32_166 ();
 DECAPx1_ASAP7_75t_SL FILLER_32_188 ();
 FILLERxp5_ASAP7_75t_SL FILLER_32_192 ();
 DECAPx10_ASAP7_75t_SL FILLER_32_196 ();
 DECAPx10_ASAP7_75t_SL FILLER_32_218 ();
 DECAPx10_ASAP7_75t_SL FILLER_32_240 ();
 DECAPx6_ASAP7_75t_SL FILLER_32_262 ();
 DECAPx2_ASAP7_75t_SL FILLER_32_276 ();
 FILLERxp5_ASAP7_75t_SL FILLER_32_282 ();
 DECAPx1_ASAP7_75t_SL FILLER_33_2 ();
 FILLERxp5_ASAP7_75t_SL FILLER_33_6 ();
 DECAPx2_ASAP7_75t_SL FILLER_33_12 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_33_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_33_33 ();
 DECAPx10_ASAP7_75t_SL FILLER_33_55 ();
 DECAPx10_ASAP7_75t_SL FILLER_33_77 ();
 DECAPx10_ASAP7_75t_SL FILLER_33_99 ();
 DECAPx10_ASAP7_75t_SL FILLER_33_121 ();
 DECAPx10_ASAP7_75t_SL FILLER_33_143 ();
 DECAPx6_ASAP7_75t_SL FILLER_33_165 ();
 DECAPx2_ASAP7_75t_SL FILLER_33_179 ();
 FILLERxp5_ASAP7_75t_SL FILLER_33_185 ();
 DECAPx6_ASAP7_75t_SL FILLER_33_192 ();
 DECAPx10_ASAP7_75t_SL FILLER_33_212 ();
 DECAPx10_ASAP7_75t_SL FILLER_33_234 ();
 DECAPx10_ASAP7_75t_SL FILLER_33_256 ();
 DECAPx1_ASAP7_75t_SL FILLER_33_278 ();
 FILLERxp5_ASAP7_75t_SL FILLER_33_282 ();
 DECAPx2_ASAP7_75t_SL FILLER_34_2 ();
 FILLERxp5_ASAP7_75t_SL FILLER_34_8 ();
 DECAPx1_ASAP7_75t_SL FILLER_34_12 ();
 FILLERxp5_ASAP7_75t_SL FILLER_34_16 ();
 FILLER_ASAP7_75t_SL FILLER_34_23 ();
 DECAPx4_ASAP7_75t_SL FILLER_34_28 ();
 FILLER_ASAP7_75t_SL FILLER_34_38 ();
 DECAPx10_ASAP7_75t_SL FILLER_34_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_34_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_34_90 ();
 FILLER_ASAP7_75t_SL FILLER_34_115 ();
 FILLER_ASAP7_75t_SL FILLER_34_123 ();
 DECAPx6_ASAP7_75t_SL FILLER_34_131 ();
 FILLERxp5_ASAP7_75t_SL FILLER_34_145 ();
 DECAPx6_ASAP7_75t_SL FILLER_34_152 ();
 FILLER_ASAP7_75t_SL FILLER_34_166 ();
 DECAPx4_ASAP7_75t_SL FILLER_34_174 ();
 FILLER_ASAP7_75t_SL FILLER_34_184 ();
 FILLER_ASAP7_75t_SL FILLER_34_206 ();
 DECAPx10_ASAP7_75t_SL FILLER_34_214 ();
 DECAPx10_ASAP7_75t_SL FILLER_34_236 ();
 DECAPx10_ASAP7_75t_SL FILLER_34_258 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_34_280 ();
 DECAPx2_ASAP7_75t_SL FILLER_35_2 ();
 FILLER_ASAP7_75t_SL FILLER_35_8 ();
 DECAPx1_ASAP7_75t_SL FILLER_35_16 ();
 FILLERxp5_ASAP7_75t_SL FILLER_35_20 ();
 DECAPx2_ASAP7_75t_SL FILLER_35_27 ();
 FILLER_ASAP7_75t_SL FILLER_35_33 ();
 DECAPx10_ASAP7_75t_SL FILLER_35_41 ();
 DECAPx10_ASAP7_75t_SL FILLER_35_63 ();
 DECAPx10_ASAP7_75t_SL FILLER_35_85 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_35_107 ();
 DECAPx6_ASAP7_75t_SL FILLER_35_130 ();
 FILLERxp5_ASAP7_75t_SL FILLER_35_144 ();
 FILLER_ASAP7_75t_SL FILLER_35_151 ();
 DECAPx4_ASAP7_75t_SL FILLER_35_159 ();
 FILLERxp5_ASAP7_75t_SL FILLER_35_169 ();
 FILLER_ASAP7_75t_SL FILLER_35_176 ();
 DECAPx1_ASAP7_75t_SL FILLER_35_184 ();
 FILLERxp5_ASAP7_75t_SL FILLER_35_188 ();
 DECAPx2_ASAP7_75t_SL FILLER_35_195 ();
 FILLER_ASAP7_75t_SL FILLER_35_204 ();
 DECAPx10_ASAP7_75t_SL FILLER_35_212 ();
 DECAPx6_ASAP7_75t_SL FILLER_35_234 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_35_248 ();
 DECAPx10_ASAP7_75t_SL FILLER_35_256 ();
 DECAPx1_ASAP7_75t_SL FILLER_35_278 ();
 FILLERxp5_ASAP7_75t_SL FILLER_35_282 ();
 FILLER_ASAP7_75t_SL FILLER_36_2 ();
 FILLER_ASAP7_75t_SL FILLER_36_9 ();
 DECAPx10_ASAP7_75t_SL FILLER_36_31 ();
 DECAPx10_ASAP7_75t_SL FILLER_36_53 ();
 DECAPx10_ASAP7_75t_SL FILLER_36_75 ();
 DECAPx2_ASAP7_75t_SL FILLER_36_97 ();
 FILLERxp5_ASAP7_75t_SL FILLER_36_103 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_36_124 ();
 DECAPx1_ASAP7_75t_SL FILLER_36_133 ();
 DECAPx1_ASAP7_75t_SL FILLER_36_157 ();
 DECAPx1_ASAP7_75t_SL FILLER_36_181 ();
 FILLERxp5_ASAP7_75t_SL FILLER_36_185 ();
 FILLER_ASAP7_75t_SL FILLER_36_206 ();
 DECAPx10_ASAP7_75t_SL FILLER_36_214 ();
 DECAPx6_ASAP7_75t_SL FILLER_36_236 ();
 FILLERxp5_ASAP7_75t_SL FILLER_36_250 ();
 DECAPx10_ASAP7_75t_SL FILLER_36_256 ();
 DECAPx1_ASAP7_75t_SL FILLER_36_278 ();
 FILLERxp5_ASAP7_75t_SL FILLER_36_282 ();
 FILLER_ASAP7_75t_SL FILLER_37_2 ();
 FILLER_ASAP7_75t_SL FILLER_37_7 ();
 DECAPx1_ASAP7_75t_SL FILLER_37_29 ();
 FILLERxp5_ASAP7_75t_SL FILLER_37_33 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_40 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_62 ();
 DECAPx6_ASAP7_75t_SL FILLER_37_84 ();
 DECAPx2_ASAP7_75t_SL FILLER_37_98 ();
 FILLER_ASAP7_75t_SL FILLER_37_107 ();
 FILLER_ASAP7_75t_SL FILLER_37_115 ();
 DECAPx2_ASAP7_75t_SL FILLER_37_123 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_37_129 ();
 DECAPx2_ASAP7_75t_SL FILLER_37_152 ();
 FILLER_ASAP7_75t_SL FILLER_37_178 ();
 FILLER_ASAP7_75t_SL FILLER_37_186 ();
 DECAPx4_ASAP7_75t_SL FILLER_37_191 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_37_201 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_207 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_229 ();
 DECAPx10_ASAP7_75t_SL FILLER_37_251 ();
 DECAPx4_ASAP7_75t_SL FILLER_37_273 ();
 FILLER_ASAP7_75t_SL FILLER_38_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_38_26 ();
 DECAPx10_ASAP7_75t_SL FILLER_38_48 ();
 DECAPx10_ASAP7_75t_SL FILLER_38_70 ();
 DECAPx10_ASAP7_75t_SL FILLER_38_92 ();
 DECAPx4_ASAP7_75t_SL FILLER_38_114 ();
 DECAPx1_ASAP7_75t_SL FILLER_38_130 ();
 FILLER_ASAP7_75t_SL FILLER_38_140 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_38_148 ();
 FILLER_ASAP7_75t_SL FILLER_38_157 ();
 DECAPx1_ASAP7_75t_SL FILLER_38_162 ();
 FILLERxp5_ASAP7_75t_SL FILLER_38_166 ();
 FILLER_ASAP7_75t_SL FILLER_38_173 ();
 DECAPx10_ASAP7_75t_SL FILLER_38_181 ();
 DECAPx10_ASAP7_75t_SL FILLER_38_203 ();
 DECAPx10_ASAP7_75t_SL FILLER_38_225 ();
 DECAPx10_ASAP7_75t_SL FILLER_38_247 ();
 DECAPx6_ASAP7_75t_SL FILLER_38_269 ();
 DECAPx2_ASAP7_75t_SL FILLER_39_2 ();
 FILLER_ASAP7_75t_SL FILLER_39_8 ();
 FILLER_ASAP7_75t_SL FILLER_39_16 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_21 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_43 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_65 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_87 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_109 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_39_131 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_137 ();
 FILLERxp5_ASAP7_75t_SL FILLER_39_159 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_163 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_185 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_207 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_229 ();
 DECAPx10_ASAP7_75t_SL FILLER_39_251 ();
 DECAPx4_ASAP7_75t_SL FILLER_39_273 ();
 FILLER_ASAP7_75t_SL FILLER_40_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_9 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_31 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_53 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_75 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_97 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_119 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_141 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_163 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_185 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_207 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_229 ();
 DECAPx10_ASAP7_75t_SL FILLER_40_251 ();
 DECAPx4_ASAP7_75t_SL FILLER_40_273 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_41_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_41_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_41_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_42_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_42_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_42_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_43_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_43_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_43_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_44_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_44_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_44_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_45_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_45_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_45_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_46_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_46_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_46_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_47_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_47_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_47_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_48_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_48_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_48_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_49_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_49_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_49_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_50_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_50_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_50_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_51_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_51_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_51_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_52_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_52_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_52_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_112 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_156 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_178 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_200 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_222 ();
 DECAPx10_ASAP7_75t_SL FILLER_53_244 ();
 DECAPx6_ASAP7_75t_SL FILLER_53_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_53_280 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_117 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_139 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_161 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_183 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_205 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_227 ();
 DECAPx10_ASAP7_75t_SL FILLER_54_249 ();
 DECAPx4_ASAP7_75t_SL FILLER_54_271 ();
 FILLER_ASAP7_75t_SL FILLER_54_281 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_90 ();
 DECAPx4_ASAP7_75t_SL FILLER_55_112 ();
 DECAPx2_ASAP7_75t_SL FILLER_55_127 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_55_133 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_55_141 ();
 DECAPx6_ASAP7_75t_SL FILLER_55_149 ();
 DECAPx1_ASAP7_75t_SL FILLER_55_163 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_55_172 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_180 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_202 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_224 ();
 DECAPx10_ASAP7_75t_SL FILLER_55_246 ();
 DECAPx6_ASAP7_75t_SL FILLER_55_268 ();
 FILLERxp5_ASAP7_75t_SL FILLER_55_282 ();
endmodule
