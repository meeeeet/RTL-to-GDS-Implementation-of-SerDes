module serializer (clock,
    dout,
    enable,
    din);
 input clock;
 output dout;
 input enable;
 input [15:0] din;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire clknet_0_clock;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire net4;
 wire net3;
 wire _064_;
 wire _065_;
 wire net2;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire net1;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire clknet_1_0__leaf_clock;
 wire clknet_1_1__leaf_clock;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;

 TAPCELL_ASAP7_75t_R PHY_5 ();
 TAPCELL_ASAP7_75t_R PHY_4 ();
 INVx1_ASAP7_75t_R _101_ (.A(_014_),
    .Y(_064_));
 NAND2x1_ASAP7_75t_R _102_ (.A(net29),
    .B(_018_),
    .Y(_065_));
 TAPCELL_ASAP7_75t_R PHY_3 ();
 OA211x2_ASAP7_75t_R _104_ (.A1(net29),
    .A2(_064_),
    .B(_065_),
    .C(net27),
    .Y(_067_));
 INVx1_ASAP7_75t_R _105_ (.A(_012_),
    .Y(_068_));
 NAND2x1_ASAP7_75t_R _106_ (.A(net29),
    .B(_016_),
    .Y(_069_));
 INVx2_ASAP7_75t_R _107_ (.A(net27),
    .Y(_070_));
 OA211x2_ASAP7_75t_R _108_ (.A1(net29),
    .A2(_068_),
    .B(_069_),
    .C(_070_),
    .Y(_071_));
 OR3x1_ASAP7_75t_R _109_ (.A(net30),
    .B(_067_),
    .C(_071_),
    .Y(_072_));
 INVx1_ASAP7_75t_R _110_ (.A(net30),
    .Y(_073_));
 INVx1_ASAP7_75t_R _111_ (.A(_015_),
    .Y(_074_));
 NAND2x1_ASAP7_75t_R _112_ (.A(net29),
    .B(_019_),
    .Y(_075_));
 OA211x2_ASAP7_75t_R _113_ (.A1(net29),
    .A2(_074_),
    .B(_075_),
    .C(net27),
    .Y(_076_));
 INVx1_ASAP7_75t_R _114_ (.A(_013_),
    .Y(_077_));
 NAND2x1_ASAP7_75t_R _115_ (.A(net29),
    .B(_017_),
    .Y(_078_));
 OA211x2_ASAP7_75t_R _116_ (.A1(net29),
    .A2(_077_),
    .B(_078_),
    .C(_070_),
    .Y(_079_));
 OR3x1_ASAP7_75t_R _117_ (.A(_073_),
    .B(_076_),
    .C(_079_),
    .Y(_080_));
 INVx1_ASAP7_75t_R _118_ (.A(_008_),
    .Y(_081_));
 NAND2x1_ASAP7_75t_R _119_ (.A(_003_),
    .B(_010_),
    .Y(_082_));
 OA211x2_ASAP7_75t_R _120_ (.A1(_003_),
    .A2(_081_),
    .B(_082_),
    .C(_000_),
    .Y(_083_));
 INVx1_ASAP7_75t_R _121_ (.A(_004_),
    .Y(_084_));
 NAND2x1_ASAP7_75t_R _122_ (.A(_003_),
    .B(_006_),
    .Y(_085_));
 INVx1_ASAP7_75t_R _123_ (.A(_000_),
    .Y(_086_));
 OA211x2_ASAP7_75t_R _124_ (.A1(_003_),
    .A2(_084_),
    .B(_085_),
    .C(_086_),
    .Y(_087_));
 OR3x1_ASAP7_75t_R _125_ (.A(_001_),
    .B(_083_),
    .C(_087_),
    .Y(_088_));
 AND2x2_ASAP7_75t_R _126_ (.A(_003_),
    .B(_011_),
    .Y(_089_));
 AO21x1_ASAP7_75t_R _127_ (.A1(_070_),
    .A2(_009_),
    .B(_089_),
    .Y(_090_));
 AND2x2_ASAP7_75t_R _128_ (.A(_001_),
    .B(_000_),
    .Y(_091_));
 AND2x2_ASAP7_75t_R _129_ (.A(_001_),
    .B(_086_),
    .Y(_092_));
 AND2x2_ASAP7_75t_R _130_ (.A(_003_),
    .B(_007_),
    .Y(_093_));
 AO21x1_ASAP7_75t_R _131_ (.A1(_070_),
    .A2(_005_),
    .B(_093_),
    .Y(_094_));
 AOI221x1_ASAP7_75t_R _132_ (.A1(_090_),
    .A2(_091_),
    .B1(_092_),
    .B2(_094_),
    .C(_002_),
    .Y(_095_));
 AO32x1_ASAP7_75t_R _133_ (.A1(_002_),
    .A2(_072_),
    .A3(_080_),
    .B1(_088_),
    .B2(_095_),
    .Y(net18));
 BUFx4_ASAP7_75t_R clkbuf_0_clock (.A(clock),
    .Y(clknet_0_clock));
 AND4x2_ASAP7_75t_R _135_ (.A(_001_),
    .B(_003_),
    .C(_000_),
    .D(_002_),
    .Y(_096_));
 TAPCELL_ASAP7_75t_R PHY_2 ();
 TAPCELL_ASAP7_75t_R PHY_1 ();
 NOR2x1_ASAP7_75t_R _138_ (.A(_019_),
    .B(net24),
    .Y(_041_));
 AO21x1_ASAP7_75t_R _139_ (.A1(net1),
    .A2(net23),
    .B(_041_),
    .Y(_021_));
 NOR2x1_ASAP7_75t_R _140_ (.A(_018_),
    .B(net24),
    .Y(_042_));
 AO21x1_ASAP7_75t_R _141_ (.A1(net8),
    .A2(net23),
    .B(_042_),
    .Y(_022_));
 NOR2x1_ASAP7_75t_R _142_ (.A(_017_),
    .B(net26),
    .Y(_043_));
 AO21x1_ASAP7_75t_R _143_ (.A1(net9),
    .A2(net23),
    .B(_043_),
    .Y(_023_));
 NOR2x1_ASAP7_75t_R _144_ (.A(_016_),
    .B(net26),
    .Y(_044_));
 AO21x1_ASAP7_75t_R _145_ (.A1(net10),
    .A2(net23),
    .B(_044_),
    .Y(_024_));
 TAPCELL_ASAP7_75t_R PHY_0 ();
 NOR2x1_ASAP7_75t_R _147_ (.A(_015_),
    .B(net24),
    .Y(_046_));
 AO21x1_ASAP7_75t_R _148_ (.A1(net11),
    .A2(net23),
    .B(_046_),
    .Y(_025_));
 NOR2x1_ASAP7_75t_R _149_ (.A(_014_),
    .B(net24),
    .Y(_047_));
 AO21x1_ASAP7_75t_R _150_ (.A1(net12),
    .A2(net23),
    .B(_047_),
    .Y(_026_));
 NOR2x1_ASAP7_75t_R _151_ (.A(_013_),
    .B(net26),
    .Y(_048_));
 AO21x1_ASAP7_75t_R _152_ (.A1(net13),
    .A2(net23),
    .B(_048_),
    .Y(_027_));
 NOR2x1_ASAP7_75t_R _153_ (.A(_012_),
    .B(net24),
    .Y(_049_));
 AO21x1_ASAP7_75t_R _154_ (.A1(net14),
    .A2(net23),
    .B(_049_),
    .Y(_028_));
 NOR2x1_ASAP7_75t_R _155_ (.A(_011_),
    .B(net26),
    .Y(_050_));
 AO21x1_ASAP7_75t_R _156_ (.A1(net15),
    .A2(net23),
    .B(_050_),
    .Y(_029_));
 NOR2x1_ASAP7_75t_R _157_ (.A(_010_),
    .B(net25),
    .Y(_051_));
 AO21x1_ASAP7_75t_R _158_ (.A1(net16),
    .A2(net23),
    .B(_051_),
    .Y(_030_));
 NOR2x1_ASAP7_75t_R _159_ (.A(_009_),
    .B(net26),
    .Y(_052_));
 AO21x1_ASAP7_75t_R _160_ (.A1(net2),
    .A2(net23),
    .B(_052_),
    .Y(_031_));
 NOR2x1_ASAP7_75t_R _161_ (.A(_008_),
    .B(net25),
    .Y(_053_));
 AO21x1_ASAP7_75t_R _162_ (.A1(net3),
    .A2(net23),
    .B(_053_),
    .Y(_032_));
 NOR2x1_ASAP7_75t_R _163_ (.A(_007_),
    .B(net26),
    .Y(_054_));
 AO21x1_ASAP7_75t_R _164_ (.A1(net4),
    .A2(net23),
    .B(_054_),
    .Y(_033_));
 NOR2x1_ASAP7_75t_R _165_ (.A(_006_),
    .B(net25),
    .Y(_055_));
 AO21x1_ASAP7_75t_R _166_ (.A1(net5),
    .A2(net23),
    .B(_055_),
    .Y(_034_));
 NOR2x1_ASAP7_75t_R _167_ (.A(_005_),
    .B(net26),
    .Y(_056_));
 AO21x1_ASAP7_75t_R _168_ (.A1(net6),
    .A2(net23),
    .B(_056_),
    .Y(_035_));
 NOR2x1_ASAP7_75t_R _169_ (.A(_004_),
    .B(net25),
    .Y(_057_));
 AO21x1_ASAP7_75t_R _170_ (.A1(net7),
    .A2(net23),
    .B(_057_),
    .Y(_036_));
 AND2x2_ASAP7_75t_R _171_ (.A(net30),
    .B(net17),
    .Y(_037_));
 XOR2x1_ASAP7_75t_R _172_ (.A(net30),
    .Y(_058_),
    .B(net28));
 AND2x2_ASAP7_75t_R _173_ (.A(net17),
    .B(_058_),
    .Y(_038_));
 OR3x1_ASAP7_75t_R _174_ (.A(net30),
    .B(net27),
    .C(net29),
    .Y(_059_));
 AO21x1_ASAP7_75t_R _175_ (.A1(_073_),
    .A2(_070_),
    .B(_086_),
    .Y(_060_));
 AND3x1_ASAP7_75t_R _176_ (.A(net17),
    .B(_059_),
    .C(_060_),
    .Y(_039_));
 XOR2x1_ASAP7_75t_R _177_ (.A(_002_),
    .Y(_061_),
    .B(_059_));
 AND2x2_ASAP7_75t_R _178_ (.A(net17),
    .B(_061_),
    .Y(_040_));
 DFFLQNx2_ASAP7_75t_R _179_ (.QN(_019_),
    .CLK(clknet_1_0__leaf_clock),
    .D(_021_));
 DFFLQNx2_ASAP7_75t_R _180_ (.QN(_018_),
    .CLK(clknet_1_1__leaf_clock),
    .D(_022_));
 DFFLQNx2_ASAP7_75t_R _181_ (.QN(_017_),
    .CLK(clknet_1_0__leaf_clock),
    .D(_023_));
 DFFLQNx2_ASAP7_75t_R _182_ (.QN(_016_),
    .CLK(clknet_1_0__leaf_clock),
    .D(_024_));
 DFFLQNx2_ASAP7_75t_R _183_ (.QN(_015_),
    .CLK(clknet_1_0__leaf_clock),
    .D(_025_));
 DFFLQNx2_ASAP7_75t_R _184_ (.QN(_014_),
    .CLK(clknet_1_0__leaf_clock),
    .D(_026_));
 DFFLQNx2_ASAP7_75t_R _185_ (.QN(_013_),
    .CLK(clknet_1_0__leaf_clock),
    .D(_027_));
 DFFLQNx2_ASAP7_75t_R _186_ (.QN(_012_),
    .CLK(clknet_1_0__leaf_clock),
    .D(_028_));
 DFFLQNx2_ASAP7_75t_R _187_ (.QN(_011_),
    .CLK(clknet_1_1__leaf_clock),
    .D(_029_));
 DFFLQNx2_ASAP7_75t_R _188_ (.QN(_010_),
    .CLK(clknet_1_1__leaf_clock),
    .D(_030_));
 DFFLQNx2_ASAP7_75t_R _189_ (.QN(_009_),
    .CLK(clknet_1_1__leaf_clock),
    .D(_031_));
 DFFLQNx2_ASAP7_75t_R _190_ (.QN(_008_),
    .CLK(clknet_1_1__leaf_clock),
    .D(_032_));
 DFFLQNx2_ASAP7_75t_R _191_ (.QN(_007_),
    .CLK(clknet_1_1__leaf_clock),
    .D(_033_));
 DFFLQNx2_ASAP7_75t_R _192_ (.QN(_006_),
    .CLK(clknet_1_1__leaf_clock),
    .D(_034_));
 DFFLQNx2_ASAP7_75t_R _193_ (.QN(_005_),
    .CLK(clknet_1_1__leaf_clock),
    .D(_035_));
 DFFLQNx2_ASAP7_75t_R _194_ (.QN(_004_),
    .CLK(clknet_1_1__leaf_clock),
    .D(_036_));
 DFFLQNx2_ASAP7_75t_R _195_ (.QN(_001_),
    .CLK(net22),
    .D(_037_));
 DFFLQNx2_ASAP7_75t_R _196_ (.QN(_003_),
    .CLK(net21),
    .D(_038_));
 DFFLQNx2_ASAP7_75t_R _197_ (.QN(_000_),
    .CLK(net20),
    .D(_039_));
 DFFLQNx2_ASAP7_75t_R _198_ (.QN(_002_),
    .CLK(net19),
    .D(_040_));
 TAPCELL_ASAP7_75t_R PHY_6 ();
 TAPCELL_ASAP7_75t_R PHY_7 ();
 TAPCELL_ASAP7_75t_R PHY_8 ();
 TAPCELL_ASAP7_75t_R PHY_9 ();
 TAPCELL_ASAP7_75t_R PHY_10 ();
 TAPCELL_ASAP7_75t_R PHY_11 ();
 TAPCELL_ASAP7_75t_R PHY_12 ();
 TAPCELL_ASAP7_75t_R PHY_13 ();
 TAPCELL_ASAP7_75t_R PHY_14 ();
 TAPCELL_ASAP7_75t_R PHY_15 ();
 TAPCELL_ASAP7_75t_R PHY_16 ();
 TAPCELL_ASAP7_75t_R PHY_17 ();
 TAPCELL_ASAP7_75t_R PHY_18 ();
 TAPCELL_ASAP7_75t_R PHY_19 ();
 TAPCELL_ASAP7_75t_R PHY_20 ();
 TAPCELL_ASAP7_75t_R PHY_21 ();
 TAPCELL_ASAP7_75t_R PHY_22 ();
 TAPCELL_ASAP7_75t_R PHY_23 ();
 TAPCELL_ASAP7_75t_R PHY_24 ();
 TAPCELL_ASAP7_75t_R PHY_25 ();
 TAPCELL_ASAP7_75t_R PHY_26 ();
 TAPCELL_ASAP7_75t_R PHY_27 ();
 TAPCELL_ASAP7_75t_R PHY_28 ();
 TAPCELL_ASAP7_75t_R PHY_29 ();
 TAPCELL_ASAP7_75t_R PHY_30 ();
 TAPCELL_ASAP7_75t_R PHY_31 ();
 TAPCELL_ASAP7_75t_R PHY_32 ();
 TAPCELL_ASAP7_75t_R PHY_33 ();
 TAPCELL_ASAP7_75t_R PHY_34 ();
 TAPCELL_ASAP7_75t_R PHY_35 ();
 TAPCELL_ASAP7_75t_R PHY_36 ();
 TAPCELL_ASAP7_75t_R PHY_37 ();
 TAPCELL_ASAP7_75t_R PHY_38 ();
 TAPCELL_ASAP7_75t_R PHY_39 ();
 TAPCELL_ASAP7_75t_R PHY_40 ();
 TAPCELL_ASAP7_75t_R PHY_41 ();
 TAPCELL_ASAP7_75t_R PHY_42 ();
 TAPCELL_ASAP7_75t_R PHY_43 ();
 TAPCELL_ASAP7_75t_R PHY_44 ();
 TAPCELL_ASAP7_75t_R PHY_45 ();
 TAPCELL_ASAP7_75t_R PHY_46 ();
 TAPCELL_ASAP7_75t_R PHY_47 ();
 TAPCELL_ASAP7_75t_R PHY_48 ();
 TAPCELL_ASAP7_75t_R PHY_49 ();
 TAPCELL_ASAP7_75t_R PHY_50 ();
 TAPCELL_ASAP7_75t_R PHY_51 ();
 TAPCELL_ASAP7_75t_R PHY_52 ();
 TAPCELL_ASAP7_75t_R PHY_53 ();
 TAPCELL_ASAP7_75t_R PHY_54 ();
 TAPCELL_ASAP7_75t_R PHY_55 ();
 TAPCELL_ASAP7_75t_R PHY_56 ();
 TAPCELL_ASAP7_75t_R PHY_57 ();
 TAPCELL_ASAP7_75t_R PHY_58 ();
 TAPCELL_ASAP7_75t_R PHY_59 ();
 TAPCELL_ASAP7_75t_R PHY_60 ();
 TAPCELL_ASAP7_75t_R PHY_61 ();
 TAPCELL_ASAP7_75t_R PHY_62 ();
 TAPCELL_ASAP7_75t_R PHY_63 ();
 TAPCELL_ASAP7_75t_R PHY_64 ();
 TAPCELL_ASAP7_75t_R PHY_65 ();
 TAPCELL_ASAP7_75t_R PHY_66 ();
 TAPCELL_ASAP7_75t_R PHY_67 ();
 TAPCELL_ASAP7_75t_R PHY_68 ();
 TAPCELL_ASAP7_75t_R PHY_69 ();
 TAPCELL_ASAP7_75t_R PHY_70 ();
 TAPCELL_ASAP7_75t_R PHY_71 ();
 TAPCELL_ASAP7_75t_R PHY_72 ();
 TAPCELL_ASAP7_75t_R PHY_73 ();
 TAPCELL_ASAP7_75t_R PHY_74 ();
 TAPCELL_ASAP7_75t_R PHY_75 ();
 TAPCELL_ASAP7_75t_R PHY_76 ();
 TAPCELL_ASAP7_75t_R PHY_77 ();
 TAPCELL_ASAP7_75t_R PHY_78 ();
 TAPCELL_ASAP7_75t_R PHY_79 ();
 TAPCELL_ASAP7_75t_R PHY_80 ();
 TAPCELL_ASAP7_75t_R PHY_81 ();
 TAPCELL_ASAP7_75t_R PHY_82 ();
 TAPCELL_ASAP7_75t_R PHY_83 ();
 BUFx2_ASAP7_75t_R input1 (.A(din[0]),
    .Y(net1));
 BUFx2_ASAP7_75t_R input2 (.A(din[10]),
    .Y(net2));
 BUFx2_ASAP7_75t_R input3 (.A(din[11]),
    .Y(net3));
 BUFx2_ASAP7_75t_R input4 (.A(din[12]),
    .Y(net4));
 BUFx2_ASAP7_75t_R input5 (.A(din[13]),
    .Y(net5));
 BUFx2_ASAP7_75t_R input6 (.A(din[14]),
    .Y(net6));
 BUFx2_ASAP7_75t_R input7 (.A(din[15]),
    .Y(net7));
 BUFx2_ASAP7_75t_R input8 (.A(din[1]),
    .Y(net8));
 BUFx2_ASAP7_75t_R input9 (.A(din[2]),
    .Y(net9));
 BUFx2_ASAP7_75t_R input10 (.A(din[3]),
    .Y(net10));
 BUFx2_ASAP7_75t_R input11 (.A(din[4]),
    .Y(net11));
 BUFx2_ASAP7_75t_R input12 (.A(din[5]),
    .Y(net12));
 BUFx2_ASAP7_75t_R input13 (.A(din[6]),
    .Y(net13));
 BUFx2_ASAP7_75t_R input14 (.A(din[7]),
    .Y(net14));
 BUFx2_ASAP7_75t_R input15 (.A(din[8]),
    .Y(net15));
 BUFx2_ASAP7_75t_R input16 (.A(din[9]),
    .Y(net16));
 BUFx2_ASAP7_75t_R input17 (.A(enable),
    .Y(net17));
 BUFx2_ASAP7_75t_R output18 (.A(net18),
    .Y(dout));
 INVx1_ASAP7_75t_R _134__1 (.A(clknet_1_1__leaf_clock),
    .Y(net19));
 INVx1_ASAP7_75t_R _134__2 (.A(clknet_1_0__leaf_clock),
    .Y(net20));
 INVx1_ASAP7_75t_R _134__3 (.A(clknet_1_1__leaf_clock),
    .Y(net21));
 INVx1_ASAP7_75t_R _134__4 (.A(clknet_1_1__leaf_clock),
    .Y(net22));
 BUFx4_ASAP7_75t_R clkbuf_1_0__f_clock (.A(clknet_0_clock),
    .Y(clknet_1_0__leaf_clock));
 BUFx4_ASAP7_75t_R clkbuf_1_1__f_clock (.A(clknet_0_clock),
    .Y(clknet_1_1__leaf_clock));
 BUFx6f_ASAP7_75t_R split5 (.A(_096_),
    .Y(net23));
 BUFx6f_ASAP7_75t_R rebuffer6 (.A(_096_),
    .Y(net24));
 BUFx3_ASAP7_75t_R rebuffer7 (.A(_096_),
    .Y(net25));
 BUFx6f_ASAP7_75t_R rebuffer8 (.A(_096_),
    .Y(net26));
 BUFx3_ASAP7_75t_R rebuffer9 (.A(_003_),
    .Y(net27));
 BUFx2_ASAP7_75t_R rebuffer10 (.A(net27),
    .Y(net28));
 BUFx3_ASAP7_75t_R rebuffer11 (.A(_000_),
    .Y(net29));
 BUFx2_ASAP7_75t_R rebuffer12 (.A(_001_),
    .Y(net30));
 DECAPx10_ASAP7_75t_R FILLER_0_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82 ();
 DECAPx4_ASAP7_75t_R FILLER_0_88 ();
 FILLER_ASAP7_75t_R FILLER_0_98 ();
 DECAPx6_ASAP7_75t_R FILLER_0_105 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_0_119 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149 ();
 DECAPx10_ASAP7_75t_R FILLER_0_171 ();
 DECAPx6_ASAP7_75t_R FILLER_0_193 ();
 DECAPx1_ASAP7_75t_R FILLER_0_207 ();
 DECAPx10_ASAP7_75t_R FILLER_1_2 ();
 DECAPx10_ASAP7_75t_R FILLER_1_24 ();
 DECAPx10_ASAP7_75t_R FILLER_1_46 ();
 DECAPx10_ASAP7_75t_R FILLER_1_68 ();
 DECAPx10_ASAP7_75t_R FILLER_1_90 ();
 DECAPx10_ASAP7_75t_R FILLER_1_112 ();
 DECAPx10_ASAP7_75t_R FILLER_1_134 ();
 DECAPx10_ASAP7_75t_R FILLER_1_156 ();
 DECAPx10_ASAP7_75t_R FILLER_1_178 ();
 DECAPx4_ASAP7_75t_R FILLER_1_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_210 ();
 DECAPx10_ASAP7_75t_R FILLER_2_2 ();
 DECAPx10_ASAP7_75t_R FILLER_2_24 ();
 DECAPx10_ASAP7_75t_R FILLER_2_46 ();
 DECAPx10_ASAP7_75t_R FILLER_2_68 ();
 DECAPx10_ASAP7_75t_R FILLER_2_90 ();
 DECAPx10_ASAP7_75t_R FILLER_2_112 ();
 DECAPx10_ASAP7_75t_R FILLER_2_134 ();
 DECAPx10_ASAP7_75t_R FILLER_2_156 ();
 DECAPx10_ASAP7_75t_R FILLER_2_178 ();
 DECAPx4_ASAP7_75t_R FILLER_2_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_210 ();
 DECAPx10_ASAP7_75t_R FILLER_3_2 ();
 DECAPx10_ASAP7_75t_R FILLER_3_24 ();
 DECAPx10_ASAP7_75t_R FILLER_3_46 ();
 DECAPx10_ASAP7_75t_R FILLER_3_68 ();
 DECAPx10_ASAP7_75t_R FILLER_3_90 ();
 DECAPx10_ASAP7_75t_R FILLER_3_112 ();
 DECAPx10_ASAP7_75t_R FILLER_3_134 ();
 DECAPx10_ASAP7_75t_R FILLER_3_156 ();
 DECAPx10_ASAP7_75t_R FILLER_3_178 ();
 DECAPx4_ASAP7_75t_R FILLER_3_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_210 ();
 DECAPx10_ASAP7_75t_R FILLER_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_4_24 ();
 DECAPx10_ASAP7_75t_R FILLER_4_46 ();
 DECAPx10_ASAP7_75t_R FILLER_4_68 ();
 DECAPx10_ASAP7_75t_R FILLER_4_90 ();
 DECAPx10_ASAP7_75t_R FILLER_4_112 ();
 DECAPx10_ASAP7_75t_R FILLER_4_134 ();
 DECAPx10_ASAP7_75t_R FILLER_4_156 ();
 DECAPx10_ASAP7_75t_R FILLER_4_178 ();
 DECAPx4_ASAP7_75t_R FILLER_4_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_210 ();
 DECAPx10_ASAP7_75t_R FILLER_5_2 ();
 DECAPx10_ASAP7_75t_R FILLER_5_24 ();
 DECAPx10_ASAP7_75t_R FILLER_5_46 ();
 DECAPx10_ASAP7_75t_R FILLER_5_68 ();
 DECAPx10_ASAP7_75t_R FILLER_5_90 ();
 DECAPx10_ASAP7_75t_R FILLER_5_112 ();
 DECAPx10_ASAP7_75t_R FILLER_5_134 ();
 DECAPx10_ASAP7_75t_R FILLER_5_156 ();
 DECAPx10_ASAP7_75t_R FILLER_5_178 ();
 DECAPx4_ASAP7_75t_R FILLER_5_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_210 ();
 DECAPx10_ASAP7_75t_R FILLER_6_2 ();
 DECAPx10_ASAP7_75t_R FILLER_6_24 ();
 DECAPx10_ASAP7_75t_R FILLER_6_46 ();
 DECAPx10_ASAP7_75t_R FILLER_6_68 ();
 DECAPx10_ASAP7_75t_R FILLER_6_90 ();
 DECAPx10_ASAP7_75t_R FILLER_6_112 ();
 DECAPx10_ASAP7_75t_R FILLER_6_134 ();
 DECAPx10_ASAP7_75t_R FILLER_6_156 ();
 DECAPx10_ASAP7_75t_R FILLER_6_178 ();
 DECAPx4_ASAP7_75t_R FILLER_6_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_210 ();
 DECAPx10_ASAP7_75t_R FILLER_7_2 ();
 DECAPx10_ASAP7_75t_R FILLER_7_24 ();
 DECAPx10_ASAP7_75t_R FILLER_7_46 ();
 DECAPx10_ASAP7_75t_R FILLER_7_68 ();
 DECAPx10_ASAP7_75t_R FILLER_7_90 ();
 DECAPx10_ASAP7_75t_R FILLER_7_112 ();
 DECAPx10_ASAP7_75t_R FILLER_7_134 ();
 DECAPx10_ASAP7_75t_R FILLER_7_156 ();
 DECAPx10_ASAP7_75t_R FILLER_7_178 ();
 DECAPx4_ASAP7_75t_R FILLER_7_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_210 ();
 DECAPx10_ASAP7_75t_R FILLER_8_2 ();
 DECAPx10_ASAP7_75t_R FILLER_8_24 ();
 DECAPx10_ASAP7_75t_R FILLER_8_46 ();
 DECAPx10_ASAP7_75t_R FILLER_8_68 ();
 DECAPx10_ASAP7_75t_R FILLER_8_90 ();
 DECAPx10_ASAP7_75t_R FILLER_8_112 ();
 DECAPx10_ASAP7_75t_R FILLER_8_134 ();
 DECAPx10_ASAP7_75t_R FILLER_8_156 ();
 DECAPx10_ASAP7_75t_R FILLER_8_178 ();
 DECAPx4_ASAP7_75t_R FILLER_8_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_210 ();
 DECAPx10_ASAP7_75t_R FILLER_9_2 ();
 DECAPx10_ASAP7_75t_R FILLER_9_24 ();
 DECAPx10_ASAP7_75t_R FILLER_9_46 ();
 DECAPx10_ASAP7_75t_R FILLER_9_68 ();
 DECAPx10_ASAP7_75t_R FILLER_9_90 ();
 DECAPx10_ASAP7_75t_R FILLER_9_112 ();
 DECAPx10_ASAP7_75t_R FILLER_9_134 ();
 DECAPx10_ASAP7_75t_R FILLER_9_156 ();
 DECAPx10_ASAP7_75t_R FILLER_9_178 ();
 DECAPx4_ASAP7_75t_R FILLER_9_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_210 ();
 DECAPx10_ASAP7_75t_R FILLER_10_2 ();
 DECAPx10_ASAP7_75t_R FILLER_10_24 ();
 DECAPx10_ASAP7_75t_R FILLER_10_46 ();
 DECAPx10_ASAP7_75t_R FILLER_10_68 ();
 DECAPx10_ASAP7_75t_R FILLER_10_90 ();
 DECAPx10_ASAP7_75t_R FILLER_10_112 ();
 DECAPx10_ASAP7_75t_R FILLER_10_134 ();
 DECAPx10_ASAP7_75t_R FILLER_10_156 ();
 DECAPx10_ASAP7_75t_R FILLER_10_178 ();
 DECAPx4_ASAP7_75t_R FILLER_10_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_210 ();
 DECAPx10_ASAP7_75t_R FILLER_11_2 ();
 DECAPx10_ASAP7_75t_R FILLER_11_24 ();
 DECAPx10_ASAP7_75t_R FILLER_11_46 ();
 DECAPx10_ASAP7_75t_R FILLER_11_68 ();
 DECAPx10_ASAP7_75t_R FILLER_11_90 ();
 DECAPx10_ASAP7_75t_R FILLER_11_112 ();
 DECAPx10_ASAP7_75t_R FILLER_11_134 ();
 DECAPx10_ASAP7_75t_R FILLER_11_156 ();
 DECAPx10_ASAP7_75t_R FILLER_11_178 ();
 DECAPx4_ASAP7_75t_R FILLER_11_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_210 ();
 DECAPx10_ASAP7_75t_R FILLER_12_2 ();
 DECAPx10_ASAP7_75t_R FILLER_12_24 ();
 DECAPx10_ASAP7_75t_R FILLER_12_46 ();
 DECAPx4_ASAP7_75t_R FILLER_12_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_12_78 ();
 DECAPx1_ASAP7_75t_R FILLER_12_102 ();
 DECAPx2_ASAP7_75t_R FILLER_12_112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_12_118 ();
 DECAPx10_ASAP7_75t_R FILLER_12_127 ();
 DECAPx10_ASAP7_75t_R FILLER_12_149 ();
 DECAPx10_ASAP7_75t_R FILLER_12_171 ();
 DECAPx6_ASAP7_75t_R FILLER_12_193 ();
 DECAPx1_ASAP7_75t_R FILLER_12_207 ();
 DECAPx2_ASAP7_75t_R FILLER_13_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_13_8 ();
 DECAPx10_ASAP7_75t_R FILLER_13_16 ();
 DECAPx10_ASAP7_75t_R FILLER_13_38 ();
 DECAPx10_ASAP7_75t_R FILLER_13_60 ();
 FILLER_ASAP7_75t_R FILLER_13_82 ();
 FILLER_ASAP7_75t_R FILLER_13_90 ();
 FILLER_ASAP7_75t_R FILLER_13_113 ();
 DECAPx10_ASAP7_75t_R FILLER_13_136 ();
 DECAPx10_ASAP7_75t_R FILLER_13_158 ();
 DECAPx10_ASAP7_75t_R FILLER_13_180 ();
 DECAPx2_ASAP7_75t_R FILLER_13_202 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_13_208 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_14_2 ();
 DECAPx10_ASAP7_75t_R FILLER_14_26 ();
 DECAPx10_ASAP7_75t_R FILLER_14_48 ();
 DECAPx6_ASAP7_75t_R FILLER_14_70 ();
 DECAPx4_ASAP7_75t_R FILLER_14_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_14_100 ();
 DECAPx4_ASAP7_75t_R FILLER_14_109 ();
 FILLER_ASAP7_75t_R FILLER_14_119 ();
 DECAPx10_ASAP7_75t_R FILLER_14_127 ();
 DECAPx10_ASAP7_75t_R FILLER_14_149 ();
 DECAPx10_ASAP7_75t_R FILLER_14_171 ();
 DECAPx6_ASAP7_75t_R FILLER_14_193 ();
 DECAPx1_ASAP7_75t_R FILLER_14_207 ();
 DECAPx1_ASAP7_75t_R FILLER_15_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_6 ();
 FILLER_ASAP7_75t_R FILLER_15_13 ();
 FILLER_ASAP7_75t_R FILLER_15_21 ();
 DECAPx6_ASAP7_75t_R FILLER_15_29 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_15_43 ();
 DECAPx6_ASAP7_75t_R FILLER_15_52 ();
 DECAPx1_ASAP7_75t_R FILLER_15_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_70 ();
 DECAPx10_ASAP7_75t_R FILLER_15_75 ();
 DECAPx10_ASAP7_75t_R FILLER_15_97 ();
 DECAPx1_ASAP7_75t_R FILLER_15_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_123 ();
 DECAPx10_ASAP7_75t_R FILLER_15_130 ();
 DECAPx10_ASAP7_75t_R FILLER_15_152 ();
 DECAPx10_ASAP7_75t_R FILLER_15_174 ();
 DECAPx2_ASAP7_75t_R FILLER_15_196 ();
 FILLER_ASAP7_75t_R FILLER_15_202 ();
 FILLER_ASAP7_75t_R FILLER_15_209 ();
 FILLER_ASAP7_75t_R FILLER_16_2 ();
 DECAPx4_ASAP7_75t_R FILLER_16_9 ();
 DECAPx10_ASAP7_75t_R FILLER_16_40 ();
 DECAPx2_ASAP7_75t_R FILLER_16_62 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_16_68 ();
 DECAPx2_ASAP7_75t_R FILLER_16_92 ();
 FILLER_ASAP7_75t_R FILLER_16_98 ();
 DECAPx4_ASAP7_75t_R FILLER_16_106 ();
 FILLER_ASAP7_75t_R FILLER_16_116 ();
 DECAPx10_ASAP7_75t_R FILLER_16_139 ();
 DECAPx10_ASAP7_75t_R FILLER_16_161 ();
 DECAPx10_ASAP7_75t_R FILLER_16_183 ();
 DECAPx2_ASAP7_75t_R FILLER_16_205 ();
 DECAPx10_ASAP7_75t_R FILLER_17_2 ();
 FILLER_ASAP7_75t_R FILLER_17_24 ();
 DECAPx4_ASAP7_75t_R FILLER_17_29 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_17_39 ();
 DECAPx4_ASAP7_75t_R FILLER_17_48 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_17_58 ();
 FILLER_ASAP7_75t_R FILLER_17_64 ();
 DECAPx2_ASAP7_75t_R FILLER_17_71 ();
 DECAPx1_ASAP7_75t_R FILLER_17_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_102 ();
 FILLER_ASAP7_75t_R FILLER_17_109 ();
 DECAPx2_ASAP7_75t_R FILLER_17_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_123 ();
 DECAPx10_ASAP7_75t_R FILLER_17_130 ();
 DECAPx10_ASAP7_75t_R FILLER_17_152 ();
 DECAPx10_ASAP7_75t_R FILLER_17_174 ();
 DECAPx6_ASAP7_75t_R FILLER_17_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_210 ();
 DECAPx1_ASAP7_75t_R FILLER_18_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_6 ();
 DECAPx2_ASAP7_75t_R FILLER_18_12 ();
 FILLER_ASAP7_75t_R FILLER_18_18 ();
 FILLER_ASAP7_75t_R FILLER_18_26 ();
 FILLER_ASAP7_75t_R FILLER_18_34 ();
 FILLER_ASAP7_75t_R FILLER_18_43 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_18_53 ();
 DECAPx2_ASAP7_75t_R FILLER_18_68 ();
 FILLER_ASAP7_75t_R FILLER_18_81 ();
 FILLER_ASAP7_75t_R FILLER_18_89 ();
 DECAPx1_ASAP7_75t_R FILLER_18_97 ();
 DECAPx1_ASAP7_75t_R FILLER_18_107 ();
 DECAPx10_ASAP7_75t_R FILLER_18_117 ();
 DECAPx10_ASAP7_75t_R FILLER_18_139 ();
 DECAPx10_ASAP7_75t_R FILLER_18_161 ();
 DECAPx10_ASAP7_75t_R FILLER_18_183 ();
 DECAPx2_ASAP7_75t_R FILLER_18_205 ();
 DECAPx4_ASAP7_75t_R FILLER_19_2 ();
 FILLER_ASAP7_75t_R FILLER_19_18 ();
 FILLER_ASAP7_75t_R FILLER_19_41 ();
 DECAPx4_ASAP7_75t_R FILLER_19_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_59 ();
 FILLER_ASAP7_75t_R FILLER_19_63 ();
 FILLER_ASAP7_75t_R FILLER_19_71 ();
 FILLER_ASAP7_75t_R FILLER_19_79 ();
 FILLER_ASAP7_75t_R FILLER_19_87 ();
 FILLER_ASAP7_75t_R FILLER_19_92 ();
 FILLER_ASAP7_75t_R FILLER_19_102 ();
 DECAPx10_ASAP7_75t_R FILLER_19_118 ();
 DECAPx10_ASAP7_75t_R FILLER_19_140 ();
 DECAPx6_ASAP7_75t_R FILLER_19_162 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_19_176 ();
 DECAPx10_ASAP7_75t_R FILLER_19_184 ();
 DECAPx1_ASAP7_75t_R FILLER_19_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_210 ();
 DECAPx4_ASAP7_75t_R FILLER_20_2 ();
 FILLER_ASAP7_75t_R FILLER_20_33 ();
 DECAPx2_ASAP7_75t_R FILLER_20_38 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_20_52 ();
 FILLER_ASAP7_75t_R FILLER_20_61 ();
 DECAPx1_ASAP7_75t_R FILLER_20_69 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_20_85 ();
 FILLER_ASAP7_75t_R FILLER_20_93 ();
 FILLER_ASAP7_75t_R FILLER_20_105 ();
 DECAPx10_ASAP7_75t_R FILLER_20_113 ();
 DECAPx10_ASAP7_75t_R FILLER_20_135 ();
 DECAPx10_ASAP7_75t_R FILLER_20_157 ();
 DECAPx10_ASAP7_75t_R FILLER_20_179 ();
 DECAPx4_ASAP7_75t_R FILLER_20_201 ();
 FILLER_ASAP7_75t_R FILLER_21_2 ();
 DECAPx4_ASAP7_75t_R FILLER_21_9 ();
 FILLER_ASAP7_75t_R FILLER_21_19 ();
 DECAPx10_ASAP7_75t_R FILLER_21_27 ();
 DECAPx1_ASAP7_75t_R FILLER_21_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_53 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_21_60 ();
 FILLER_ASAP7_75t_R FILLER_21_70 ();
 FILLER_ASAP7_75t_R FILLER_21_78 ();
 FILLER_ASAP7_75t_R FILLER_21_101 ();
 DECAPx10_ASAP7_75t_R FILLER_21_113 ();
 DECAPx10_ASAP7_75t_R FILLER_21_135 ();
 DECAPx10_ASAP7_75t_R FILLER_21_157 ();
 DECAPx6_ASAP7_75t_R FILLER_21_179 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_21_193 ();
 DECAPx4_ASAP7_75t_R FILLER_21_201 ();
 FILLER_ASAP7_75t_R FILLER_22_2 ();
 DECAPx4_ASAP7_75t_R FILLER_22_9 ();
 FILLER_ASAP7_75t_R FILLER_22_19 ();
 DECAPx6_ASAP7_75t_R FILLER_22_27 ();
 FILLER_ASAP7_75t_R FILLER_22_44 ();
 DECAPx6_ASAP7_75t_R FILLER_22_54 ();
 DECAPx1_ASAP7_75t_R FILLER_22_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_72 ();
 FILLER_ASAP7_75t_R FILLER_22_94 ();
 DECAPx1_ASAP7_75t_R FILLER_22_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_103 ();
 FILLER_ASAP7_75t_R FILLER_22_112 ();
 DECAPx10_ASAP7_75t_R FILLER_22_120 ();
 DECAPx10_ASAP7_75t_R FILLER_22_142 ();
 DECAPx10_ASAP7_75t_R FILLER_22_164 ();
 DECAPx10_ASAP7_75t_R FILLER_22_186 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_22_208 ();
 FILLER_ASAP7_75t_R FILLER_23_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_23_25 ();
 DECAPx2_ASAP7_75t_R FILLER_23_34 ();
 DECAPx10_ASAP7_75t_R FILLER_23_46 ();
 DECAPx2_ASAP7_75t_R FILLER_23_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_74 ();
 DECAPx1_ASAP7_75t_R FILLER_23_78 ();
 DECAPx2_ASAP7_75t_R FILLER_23_85 ();
 FILLER_ASAP7_75t_R FILLER_23_91 ();
 DECAPx2_ASAP7_75t_R FILLER_23_99 ();
 FILLER_ASAP7_75t_R FILLER_23_105 ();
 DECAPx10_ASAP7_75t_R FILLER_23_115 ();
 DECAPx10_ASAP7_75t_R FILLER_23_137 ();
 DECAPx10_ASAP7_75t_R FILLER_23_159 ();
 DECAPx10_ASAP7_75t_R FILLER_23_181 ();
 DECAPx2_ASAP7_75t_R FILLER_23_203 ();
 FILLER_ASAP7_75t_R FILLER_23_209 ();
 DECAPx1_ASAP7_75t_R FILLER_24_2 ();
 FILLER_ASAP7_75t_R FILLER_24_12 ();
 DECAPx2_ASAP7_75t_R FILLER_24_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_25 ();
 DECAPx10_ASAP7_75t_R FILLER_24_47 ();
 DECAPx10_ASAP7_75t_R FILLER_24_69 ();
 DECAPx2_ASAP7_75t_R FILLER_24_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_97 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_24_106 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_24_115 ();
 DECAPx10_ASAP7_75t_R FILLER_24_121 ();
 DECAPx10_ASAP7_75t_R FILLER_24_143 ();
 DECAPx10_ASAP7_75t_R FILLER_24_165 ();
 DECAPx10_ASAP7_75t_R FILLER_24_187 ();
 FILLER_ASAP7_75t_R FILLER_24_209 ();
 DECAPx4_ASAP7_75t_R FILLER_25_2 ();
 FILLER_ASAP7_75t_R FILLER_25_12 ();
 FILLER_ASAP7_75t_R FILLER_25_35 ();
 FILLER_ASAP7_75t_R FILLER_25_40 ();
 FILLER_ASAP7_75t_R FILLER_25_48 ();
 FILLER_ASAP7_75t_R FILLER_25_58 ();
 DECAPx10_ASAP7_75t_R FILLER_25_66 ();
 DECAPx2_ASAP7_75t_R FILLER_25_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_94 ();
 FILLER_ASAP7_75t_R FILLER_25_98 ();
 DECAPx1_ASAP7_75t_R FILLER_25_106 ();
 FILLER_ASAP7_75t_R FILLER_25_131 ();
 DECAPx10_ASAP7_75t_R FILLER_25_139 ();
 DECAPx10_ASAP7_75t_R FILLER_25_161 ();
 DECAPx10_ASAP7_75t_R FILLER_25_183 ();
 DECAPx2_ASAP7_75t_R FILLER_25_205 ();
 FILLER_ASAP7_75t_R FILLER_26_2 ();
 FILLER_ASAP7_75t_R FILLER_26_9 ();
 DECAPx4_ASAP7_75t_R FILLER_26_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_27 ();
 DECAPx10_ASAP7_75t_R FILLER_26_34 ();
 DECAPx2_ASAP7_75t_R FILLER_26_56 ();
 FILLER_ASAP7_75t_R FILLER_26_62 ();
 DECAPx10_ASAP7_75t_R FILLER_26_70 ();
 FILLER_ASAP7_75t_R FILLER_26_92 ();
 FILLER_ASAP7_75t_R FILLER_26_100 ();
 DECAPx10_ASAP7_75t_R FILLER_26_108 ();
 DECAPx1_ASAP7_75t_R FILLER_26_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_134 ();
 DECAPx10_ASAP7_75t_R FILLER_26_141 ();
 DECAPx10_ASAP7_75t_R FILLER_26_163 ();
 DECAPx10_ASAP7_75t_R FILLER_26_185 ();
 DECAPx1_ASAP7_75t_R FILLER_26_207 ();
 DECAPx10_ASAP7_75t_R FILLER_27_2 ();
 DECAPx10_ASAP7_75t_R FILLER_27_24 ();
 DECAPx2_ASAP7_75t_R FILLER_27_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_52 ();
 FILLER_ASAP7_75t_R FILLER_27_74 ();
 FILLER_ASAP7_75t_R FILLER_27_97 ();
 FILLER_ASAP7_75t_R FILLER_27_109 ();
 DECAPx1_ASAP7_75t_R FILLER_27_117 ();
 DECAPx10_ASAP7_75t_R FILLER_27_127 ();
 DECAPx10_ASAP7_75t_R FILLER_27_149 ();
 DECAPx10_ASAP7_75t_R FILLER_27_171 ();
 DECAPx6_ASAP7_75t_R FILLER_27_193 ();
 DECAPx1_ASAP7_75t_R FILLER_27_207 ();
 DECAPx10_ASAP7_75t_R FILLER_28_2 ();
 DECAPx10_ASAP7_75t_R FILLER_28_24 ();
 DECAPx6_ASAP7_75t_R FILLER_28_46 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_60 ();
 DECAPx4_ASAP7_75t_R FILLER_28_69 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_79 ();
 FILLER_ASAP7_75t_R FILLER_28_88 ();
 FILLER_ASAP7_75t_R FILLER_28_111 ();
 DECAPx10_ASAP7_75t_R FILLER_28_134 ();
 DECAPx10_ASAP7_75t_R FILLER_28_156 ();
 DECAPx10_ASAP7_75t_R FILLER_28_178 ();
 DECAPx4_ASAP7_75t_R FILLER_28_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_210 ();
 DECAPx10_ASAP7_75t_R FILLER_29_2 ();
 DECAPx10_ASAP7_75t_R FILLER_29_24 ();
 DECAPx10_ASAP7_75t_R FILLER_29_46 ();
 DECAPx10_ASAP7_75t_R FILLER_29_68 ();
 DECAPx4_ASAP7_75t_R FILLER_29_90 ();
 DECAPx4_ASAP7_75t_R FILLER_29_106 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_29_116 ();
 DECAPx10_ASAP7_75t_R FILLER_29_125 ();
 DECAPx10_ASAP7_75t_R FILLER_29_147 ();
 DECAPx10_ASAP7_75t_R FILLER_29_169 ();
 DECAPx6_ASAP7_75t_R FILLER_29_191 ();
 DECAPx2_ASAP7_75t_R FILLER_29_205 ();
 DECAPx10_ASAP7_75t_R FILLER_30_2 ();
 DECAPx10_ASAP7_75t_R FILLER_30_24 ();
 DECAPx10_ASAP7_75t_R FILLER_30_46 ();
 DECAPx10_ASAP7_75t_R FILLER_30_68 ();
 DECAPx10_ASAP7_75t_R FILLER_30_90 ();
 DECAPx10_ASAP7_75t_R FILLER_30_112 ();
 DECAPx10_ASAP7_75t_R FILLER_30_134 ();
 DECAPx10_ASAP7_75t_R FILLER_30_156 ();
 DECAPx10_ASAP7_75t_R FILLER_30_178 ();
 DECAPx4_ASAP7_75t_R FILLER_30_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_210 ();
 DECAPx10_ASAP7_75t_R FILLER_31_2 ();
 DECAPx10_ASAP7_75t_R FILLER_31_24 ();
 DECAPx10_ASAP7_75t_R FILLER_31_46 ();
 DECAPx10_ASAP7_75t_R FILLER_31_68 ();
 DECAPx10_ASAP7_75t_R FILLER_31_90 ();
 DECAPx10_ASAP7_75t_R FILLER_31_112 ();
 DECAPx10_ASAP7_75t_R FILLER_31_134 ();
 DECAPx10_ASAP7_75t_R FILLER_31_156 ();
 DECAPx10_ASAP7_75t_R FILLER_31_178 ();
 DECAPx4_ASAP7_75t_R FILLER_31_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_210 ();
 DECAPx10_ASAP7_75t_R FILLER_32_2 ();
 DECAPx10_ASAP7_75t_R FILLER_32_24 ();
 DECAPx10_ASAP7_75t_R FILLER_32_46 ();
 DECAPx10_ASAP7_75t_R FILLER_32_68 ();
 DECAPx10_ASAP7_75t_R FILLER_32_90 ();
 DECAPx10_ASAP7_75t_R FILLER_32_112 ();
 DECAPx10_ASAP7_75t_R FILLER_32_134 ();
 DECAPx10_ASAP7_75t_R FILLER_32_156 ();
 DECAPx10_ASAP7_75t_R FILLER_32_178 ();
 DECAPx4_ASAP7_75t_R FILLER_32_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_210 ();
 DECAPx10_ASAP7_75t_R FILLER_33_2 ();
 DECAPx10_ASAP7_75t_R FILLER_33_24 ();
 DECAPx10_ASAP7_75t_R FILLER_33_46 ();
 DECAPx10_ASAP7_75t_R FILLER_33_68 ();
 DECAPx10_ASAP7_75t_R FILLER_33_90 ();
 DECAPx10_ASAP7_75t_R FILLER_33_112 ();
 DECAPx10_ASAP7_75t_R FILLER_33_134 ();
 DECAPx10_ASAP7_75t_R FILLER_33_156 ();
 DECAPx10_ASAP7_75t_R FILLER_33_178 ();
 DECAPx4_ASAP7_75t_R FILLER_33_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_210 ();
 DECAPx10_ASAP7_75t_R FILLER_34_2 ();
 DECAPx10_ASAP7_75t_R FILLER_34_24 ();
 DECAPx10_ASAP7_75t_R FILLER_34_46 ();
 DECAPx10_ASAP7_75t_R FILLER_34_68 ();
 DECAPx10_ASAP7_75t_R FILLER_34_90 ();
 DECAPx10_ASAP7_75t_R FILLER_34_112 ();
 DECAPx10_ASAP7_75t_R FILLER_34_134 ();
 DECAPx10_ASAP7_75t_R FILLER_34_156 ();
 DECAPx10_ASAP7_75t_R FILLER_34_178 ();
 DECAPx4_ASAP7_75t_R FILLER_34_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_210 ();
 DECAPx10_ASAP7_75t_R FILLER_35_2 ();
 DECAPx10_ASAP7_75t_R FILLER_35_24 ();
 DECAPx10_ASAP7_75t_R FILLER_35_46 ();
 DECAPx10_ASAP7_75t_R FILLER_35_68 ();
 DECAPx10_ASAP7_75t_R FILLER_35_90 ();
 DECAPx10_ASAP7_75t_R FILLER_35_112 ();
 DECAPx10_ASAP7_75t_R FILLER_35_134 ();
 DECAPx10_ASAP7_75t_R FILLER_35_156 ();
 DECAPx10_ASAP7_75t_R FILLER_35_178 ();
 DECAPx4_ASAP7_75t_R FILLER_35_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_210 ();
 DECAPx10_ASAP7_75t_R FILLER_36_2 ();
 DECAPx10_ASAP7_75t_R FILLER_36_24 ();
 DECAPx10_ASAP7_75t_R FILLER_36_46 ();
 DECAPx10_ASAP7_75t_R FILLER_36_68 ();
 DECAPx10_ASAP7_75t_R FILLER_36_90 ();
 DECAPx10_ASAP7_75t_R FILLER_36_112 ();
 DECAPx10_ASAP7_75t_R FILLER_36_134 ();
 DECAPx10_ASAP7_75t_R FILLER_36_156 ();
 DECAPx10_ASAP7_75t_R FILLER_36_178 ();
 DECAPx4_ASAP7_75t_R FILLER_36_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_210 ();
 DECAPx10_ASAP7_75t_R FILLER_37_2 ();
 DECAPx10_ASAP7_75t_R FILLER_37_24 ();
 DECAPx10_ASAP7_75t_R FILLER_37_46 ();
 DECAPx10_ASAP7_75t_R FILLER_37_68 ();
 DECAPx10_ASAP7_75t_R FILLER_37_90 ();
 DECAPx10_ASAP7_75t_R FILLER_37_112 ();
 DECAPx10_ASAP7_75t_R FILLER_37_134 ();
 DECAPx10_ASAP7_75t_R FILLER_37_156 ();
 DECAPx10_ASAP7_75t_R FILLER_37_178 ();
 DECAPx4_ASAP7_75t_R FILLER_37_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_210 ();
 DECAPx10_ASAP7_75t_R FILLER_38_2 ();
 DECAPx10_ASAP7_75t_R FILLER_38_24 ();
 DECAPx10_ASAP7_75t_R FILLER_38_46 ();
 DECAPx10_ASAP7_75t_R FILLER_38_68 ();
 DECAPx10_ASAP7_75t_R FILLER_38_90 ();
 DECAPx10_ASAP7_75t_R FILLER_38_112 ();
 DECAPx10_ASAP7_75t_R FILLER_38_134 ();
 DECAPx10_ASAP7_75t_R FILLER_38_156 ();
 DECAPx10_ASAP7_75t_R FILLER_38_178 ();
 DECAPx4_ASAP7_75t_R FILLER_38_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_210 ();
 DECAPx10_ASAP7_75t_R FILLER_39_2 ();
 DECAPx10_ASAP7_75t_R FILLER_39_24 ();
 DECAPx10_ASAP7_75t_R FILLER_39_46 ();
 DECAPx10_ASAP7_75t_R FILLER_39_68 ();
 DECAPx10_ASAP7_75t_R FILLER_39_90 ();
 DECAPx10_ASAP7_75t_R FILLER_39_112 ();
 DECAPx10_ASAP7_75t_R FILLER_39_134 ();
 DECAPx10_ASAP7_75t_R FILLER_39_156 ();
 DECAPx10_ASAP7_75t_R FILLER_39_178 ();
 DECAPx4_ASAP7_75t_R FILLER_39_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_210 ();
 DECAPx10_ASAP7_75t_R FILLER_40_2 ();
 DECAPx10_ASAP7_75t_R FILLER_40_24 ();
 DECAPx10_ASAP7_75t_R FILLER_40_46 ();
 DECAPx4_ASAP7_75t_R FILLER_40_68 ();
 FILLER_ASAP7_75t_R FILLER_40_78 ();
 DECAPx10_ASAP7_75t_R FILLER_40_85 ();
 DECAPx10_ASAP7_75t_R FILLER_40_107 ();
 DECAPx10_ASAP7_75t_R FILLER_40_129 ();
 DECAPx10_ASAP7_75t_R FILLER_40_151 ();
 DECAPx10_ASAP7_75t_R FILLER_40_173 ();
 DECAPx6_ASAP7_75t_R FILLER_40_195 ();
 FILLER_ASAP7_75t_R FILLER_40_209 ();
 DECAPx10_ASAP7_75t_R FILLER_41_2 ();
 DECAPx10_ASAP7_75t_R FILLER_41_24 ();
 DECAPx6_ASAP7_75t_R FILLER_41_46 ();
 DECAPx1_ASAP7_75t_R FILLER_41_60 ();
 DECAPx10_ASAP7_75t_R FILLER_41_69 ();
 DECAPx2_ASAP7_75t_R FILLER_41_91 ();
 FILLER_ASAP7_75t_R FILLER_41_97 ();
 DECAPx6_ASAP7_75t_R FILLER_41_104 ();
 DECAPx1_ASAP7_75t_R FILLER_41_118 ();
 DECAPx2_ASAP7_75t_R FILLER_41_127 ();
 FILLER_ASAP7_75t_R FILLER_41_133 ();
 DECAPx10_ASAP7_75t_R FILLER_41_140 ();
 DECAPx10_ASAP7_75t_R FILLER_41_162 ();
 DECAPx10_ASAP7_75t_R FILLER_41_184 ();
 DECAPx1_ASAP7_75t_R FILLER_41_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_210 ();
endmodule
