// Code your design here
