module ser_top (clk,
    data_en,
    load_en,
    rst_n,
    ser_out,
    parallel_data_in);
 input clk;
 input data_en;
 input load_en;
 input rst_n;
 output ser_out;
 input [7:0] parallel_data_in;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire clknet_0_clk;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire net3;
 wire net2;
 wire _061_;
 wire net1;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire net8;
 wire net7;
 wire _118_;
 wire net6;
 wire _120_;
 wire net5;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire net4;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire \data_in_latch.data_8b_out[0] ;
 wire \data_in_latch.data_8b_out[1] ;
 wire \data_in_latch.data_8b_out[2] ;
 wire \data_in_latch.data_8b_out[3] ;
 wire \data_in_latch.data_8b_out[4] ;
 wire \data_in_latch.data_8b_out[5] ;
 wire \data_in_latch.data_8b_out[6] ;
 wire \data_in_latch.data_8b_out[7] ;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 TAPCELL_ASAP7_75t_SL PHY_9 ();
 AND2x2_ASAP7_75t_SL _133_ (.A(net11),
    .B(net3),
    .Y(_000_));
 AND2x2_ASAP7_75t_SL _134_ (.A(net11),
    .B(net4),
    .Y(_001_));
 AND2x2_ASAP7_75t_SL _135_ (.A(net11),
    .B(net5),
    .Y(_002_));
 AND2x2_ASAP7_75t_SL _136_ (.A(net11),
    .B(net6),
    .Y(_003_));
 AND2x2_ASAP7_75t_SL _137_ (.A(net11),
    .B(net7),
    .Y(_004_));
 AND2x2_ASAP7_75t_SL _138_ (.A(net11),
    .B(net8),
    .Y(_005_));
 AND2x2_ASAP7_75t_SL _139_ (.A(net11),
    .B(net9),
    .Y(_006_));
 AND2x2_ASAP7_75t_SL _140_ (.A(net11),
    .B(net10),
    .Y(_007_));
 TAPCELL_ASAP7_75t_SL PHY_8 ();
 INVx2_ASAP7_75t_SL _142_ (.A(net1),
    .Y(_118_));
 AND2x4_ASAP7_75t_SL _143_ (.A(net11),
    .B(_118_),
    .Y(_008_));
 BUFx4_ASAP7_75t_SL clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 INVx1_ASAP7_75t_SL _145_ (.A(_009_),
    .Y(net12));
 TAPCELL_ASAP7_75t_SL PHY_7 ();
 CKINVDCx5p33_ASAP7_75t_SL _147_ (.A(net2),
    .Y(_120_));
 TAPCELL_ASAP7_75t_SL PHY_6 ();
 AND3x1_ASAP7_75t_SL _149_ (.A(net11),
    .B(_120_),
    .C(_027_),
    .Y(_122_));
 INVx1_ASAP7_75t_SL _150_ (.A(net11),
    .Y(_123_));
 OA21x2_ASAP7_75t_SL _151_ (.A1(_123_),
    .A2(net2),
    .B(_009_),
    .Y(_124_));
 NOR2x1_ASAP7_75t_SL _152_ (.A(_122_),
    .B(_124_),
    .Y(_047_));
 INVx1_ASAP7_75t_SL _153_ (.A(_026_),
    .Y(_125_));
 NAND2x1_ASAP7_75t_SL _154_ (.A(net2),
    .B(_013_),
    .Y(_126_));
 TAPCELL_ASAP7_75t_SL PHY_5 ();
 OA211x2_ASAP7_75t_SL _156_ (.A1(net2),
    .A2(_125_),
    .B(_126_),
    .C(net11),
    .Y(_029_));
 INVx1_ASAP7_75t_SL _157_ (.A(_012_),
    .Y(_128_));
 NAND2x1_ASAP7_75t_SL _158_ (.A(_120_),
    .B(_025_),
    .Y(_129_));
 OA211x2_ASAP7_75t_SL _159_ (.A1(_120_),
    .A2(_128_),
    .B(_129_),
    .C(net11),
    .Y(_030_));
 INVx1_ASAP7_75t_SL _160_ (.A(_024_),
    .Y(_130_));
 NAND2x1_ASAP7_75t_SL _161_ (.A(net2),
    .B(_011_),
    .Y(_131_));
 OA211x2_ASAP7_75t_SL _162_ (.A1(net2),
    .A2(_130_),
    .B(_131_),
    .C(net11),
    .Y(_031_));
 INVx1_ASAP7_75t_SL _163_ (.A(_019_),
    .Y(_048_));
 NAND2x1_ASAP7_75t_SL _164_ (.A(_120_),
    .B(_023_),
    .Y(_049_));
 OA211x2_ASAP7_75t_SL _165_ (.A1(_120_),
    .A2(_048_),
    .B(_049_),
    .C(net11),
    .Y(_032_));
 INVx1_ASAP7_75t_SL _166_ (.A(_018_),
    .Y(_050_));
 NAND2x1_ASAP7_75t_SL _167_ (.A(_120_),
    .B(_022_),
    .Y(_051_));
 OA211x2_ASAP7_75t_SL _168_ (.A1(_120_),
    .A2(_050_),
    .B(_051_),
    .C(net11),
    .Y(_033_));
 INVx1_ASAP7_75t_SL _169_ (.A(_017_),
    .Y(_052_));
 NAND2x1_ASAP7_75t_SL _170_ (.A(_120_),
    .B(_021_),
    .Y(_053_));
 OA211x2_ASAP7_75t_SL _171_ (.A1(_120_),
    .A2(_052_),
    .B(_053_),
    .C(net11),
    .Y(_034_));
 INVx1_ASAP7_75t_SL _172_ (.A(_016_),
    .Y(_054_));
 NAND2x1_ASAP7_75t_SL _173_ (.A(_120_),
    .B(_020_),
    .Y(_055_));
 OA211x2_ASAP7_75t_SL _174_ (.A1(_120_),
    .A2(_054_),
    .B(_055_),
    .C(net11),
    .Y(_035_));
 INVx1_ASAP7_75t_SL _175_ (.A(_015_),
    .Y(_056_));
 NAND2x1_ASAP7_75t_SL _176_ (.A(_120_),
    .B(_010_),
    .Y(_057_));
 OA211x2_ASAP7_75t_SL _177_ (.A1(_120_),
    .A2(_056_),
    .B(_057_),
    .C(net11),
    .Y(_036_));
 INVx1_ASAP7_75t_SL _178_ (.A(\data_in_latch.data_8b_out[1] ),
    .Y(_058_));
 TAPCELL_ASAP7_75t_SL PHY_4 ();
 TAPCELL_ASAP7_75t_SL PHY_3 ();
 NOR2x1_ASAP7_75t_SL _181_ (.A(\data_in_latch.data_8b_out[2] ),
    .B(\data_in_latch.data_8b_out[4] ),
    .Y(_061_));
 TAPCELL_ASAP7_75t_SL PHY_2 ();
 TAPCELL_ASAP7_75t_SL PHY_1 ();
 NAND2x1_ASAP7_75t_SL _184_ (.A(\data_in_latch.data_8b_out[0] ),
    .B(\data_in_latch.data_8b_out[3] ),
    .Y(_064_));
 OR2x2_ASAP7_75t_SL _185_ (.A(\data_in_latch.data_8b_out[0] ),
    .B(\data_in_latch.data_8b_out[3] ),
    .Y(_065_));
 OA211x2_ASAP7_75t_SL _186_ (.A1(_058_),
    .A2(_061_),
    .B(_064_),
    .C(_065_),
    .Y(_066_));
 AND3x1_ASAP7_75t_SL _187_ (.A(\data_in_latch.data_8b_out[0] ),
    .B(_058_),
    .C(_061_),
    .Y(_067_));
 INVx2_ASAP7_75t_SL _188_ (.A(\data_in_latch.data_8b_out[0] ),
    .Y(_068_));
 INVx1_ASAP7_75t_SL _189_ (.A(\data_in_latch.data_8b_out[3] ),
    .Y(_069_));
 AND3x1_ASAP7_75t_SL _190_ (.A(_068_),
    .B(_069_),
    .C(\data_in_latch.data_8b_out[4] ),
    .Y(_070_));
 NOR2x1_ASAP7_75t_SL _191_ (.A(\data_in_latch.data_8b_out[0] ),
    .B(\data_in_latch.data_8b_out[3] ),
    .Y(_071_));
 TAPCELL_ASAP7_75t_SL PHY_0 ();
 AND3x1_ASAP7_75t_SL _193_ (.A(\data_in_latch.data_8b_out[0] ),
    .B(\data_in_latch.data_8b_out[1] ),
    .C(\data_in_latch.data_8b_out[3] ),
    .Y(_073_));
 OA21x2_ASAP7_75t_SL _194_ (.A1(_071_),
    .A2(_073_),
    .B(\data_in_latch.data_8b_out[2] ),
    .Y(_074_));
 OR4x1_ASAP7_75t_SL _195_ (.A(_066_),
    .B(_067_),
    .C(_070_),
    .D(_074_),
    .Y(_075_));
 NOR2x1_ASAP7_75t_SL _196_ (.A(\data_in_latch.data_8b_out[1] ),
    .B(\data_in_latch.data_8b_out[3] ),
    .Y(_076_));
 NAND2x1_ASAP7_75t_SL _197_ (.A(\data_in_latch.data_8b_out[2] ),
    .B(\data_in_latch.data_8b_out[4] ),
    .Y(_077_));
 AND2x2_ASAP7_75t_SL _198_ (.A(\data_in_latch.data_8b_out[0] ),
    .B(\data_in_latch.data_8b_out[1] ),
    .Y(_078_));
 AOI211x1_ASAP7_75t_SL _199_ (.A1(_068_),
    .A2(_076_),
    .B(_077_),
    .C(_078_),
    .Y(_079_));
 INVx1_ASAP7_75t_SL _200_ (.A(_079_),
    .Y(_080_));
 OR2x2_ASAP7_75t_SL _201_ (.A(\data_in_latch.data_8b_out[3] ),
    .B(\data_in_latch.data_8b_out[4] ),
    .Y(_081_));
 OR3x1_ASAP7_75t_SL _202_ (.A(\data_in_latch.data_8b_out[0] ),
    .B(\data_in_latch.data_8b_out[1] ),
    .C(\data_in_latch.data_8b_out[2] ),
    .Y(_082_));
 AND2x2_ASAP7_75t_SL _203_ (.A(net11),
    .B(net1),
    .Y(_083_));
 OA21x2_ASAP7_75t_SL _204_ (.A1(_081_),
    .A2(_082_),
    .B(_083_),
    .Y(_084_));
 AO32x1_ASAP7_75t_SL _205_ (.A1(_075_),
    .A2(_080_),
    .A3(_084_),
    .B1(_008_),
    .B2(_048_),
    .Y(_037_));
 INVx3_ASAP7_75t_SL _206_ (.A(\data_in_latch.data_8b_out[2] ),
    .Y(_085_));
 AND2x2_ASAP7_75t_SL _207_ (.A(\data_in_latch.data_8b_out[3] ),
    .B(\data_in_latch.data_8b_out[2] ),
    .Y(_086_));
 AO22x1_ASAP7_75t_SL _208_ (.A1(_085_),
    .A2(_071_),
    .B1(_086_),
    .B2(\data_in_latch.data_8b_out[0] ),
    .Y(_087_));
 AO21x1_ASAP7_75t_SL _209_ (.A1(\data_in_latch.data_8b_out[1] ),
    .A2(_087_),
    .B(\data_in_latch.data_8b_out[4] ),
    .Y(_088_));
 AO22x1_ASAP7_75t_SL _210_ (.A1(_050_),
    .A2(_008_),
    .B1(_083_),
    .B2(_088_),
    .Y(_038_));
 INVx1_ASAP7_75t_SL _211_ (.A(\data_in_latch.data_8b_out[4] ),
    .Y(_089_));
 AO21x1_ASAP7_75t_SL _212_ (.A1(_058_),
    .A2(_089_),
    .B(\data_in_latch.data_8b_out[3] ),
    .Y(_090_));
 NAND2x1_ASAP7_75t_SL _213_ (.A(\data_in_latch.data_8b_out[1] ),
    .B(\data_in_latch.data_8b_out[4] ),
    .Y(_091_));
 AO21x1_ASAP7_75t_SL _214_ (.A1(\data_in_latch.data_8b_out[3] ),
    .A2(_091_),
    .B(_085_),
    .Y(_092_));
 OA21x2_ASAP7_75t_SL _215_ (.A1(_068_),
    .A2(_092_),
    .B(_082_),
    .Y(_093_));
 AO32x1_ASAP7_75t_SL _216_ (.A1(_083_),
    .A2(_090_),
    .A3(_093_),
    .B1(_008_),
    .B2(_052_),
    .Y(_039_));
 MAJx2_ASAP7_75t_SL _217_ (.A(\data_in_latch.data_8b_out[0] ),
    .B(\data_in_latch.data_8b_out[3] ),
    .C(\data_in_latch.data_8b_out[4] ),
    .Y(_094_));
 NAND2x1_ASAP7_75t_SL _218_ (.A(_085_),
    .B(_094_),
    .Y(_095_));
 OA21x2_ASAP7_75t_SL _219_ (.A1(\data_in_latch.data_8b_out[4] ),
    .A2(_064_),
    .B(\data_in_latch.data_8b_out[2] ),
    .Y(_096_));
 OR4x1_ASAP7_75t_SL _220_ (.A(\data_in_latch.data_8b_out[0] ),
    .B(\data_in_latch.data_8b_out[1] ),
    .C(_085_),
    .D(_081_),
    .Y(_097_));
 OA211x2_ASAP7_75t_SL _221_ (.A1(_058_),
    .A2(_096_),
    .B(_097_),
    .C(_083_),
    .Y(_098_));
 AO32x1_ASAP7_75t_SL _222_ (.A1(net11),
    .A2(_118_),
    .A3(_054_),
    .B1(_095_),
    .B2(_098_),
    .Y(_040_));
 NAND2x1_ASAP7_75t_SL _223_ (.A(\data_in_latch.data_8b_out[2] ),
    .B(_081_),
    .Y(_099_));
 AO221x1_ASAP7_75t_SL _224_ (.A1(_085_),
    .A2(_089_),
    .B1(_099_),
    .B2(_068_),
    .C(\data_in_latch.data_8b_out[1] ),
    .Y(_100_));
 AO21x1_ASAP7_75t_SL _225_ (.A1(\data_in_latch.data_8b_out[1] ),
    .A2(_077_),
    .B(_064_),
    .Y(_101_));
 AO32x1_ASAP7_75t_SL _226_ (.A1(_083_),
    .A2(_100_),
    .A3(_101_),
    .B1(_008_),
    .B2(_056_),
    .Y(_041_));
 AO21x1_ASAP7_75t_SL _227_ (.A1(_089_),
    .A2(_086_),
    .B(_068_),
    .Y(_102_));
 AO21x1_ASAP7_75t_SL _228_ (.A1(_069_),
    .A2(\data_in_latch.data_8b_out[4] ),
    .B(_086_),
    .Y(_103_));
 AO21x1_ASAP7_75t_SL _229_ (.A1(_061_),
    .A2(_076_),
    .B(_118_),
    .Y(_104_));
 AO221x1_ASAP7_75t_SL _230_ (.A1(\data_in_latch.data_8b_out[1] ),
    .A2(_102_),
    .B1(_103_),
    .B2(_068_),
    .C(_104_),
    .Y(_105_));
 OR2x2_ASAP7_75t_SL _231_ (.A(net1),
    .B(_014_),
    .Y(_106_));
 AOI21x1_ASAP7_75t_SL _232_ (.A1(_105_),
    .A2(_106_),
    .B(_123_),
    .Y(_042_));
 NAND2x1_ASAP7_75t_SL _233_ (.A(\data_in_latch.data_8b_out[5] ),
    .B(\data_in_latch.data_8b_out[6] ),
    .Y(_107_));
 XNOR2x1_ASAP7_75t_SL _234_ (.B(_107_),
    .Y(_108_),
    .A(\data_in_latch.data_8b_out[7] ));
 NAND2x1_ASAP7_75t_SL _235_ (.A(_118_),
    .B(_013_),
    .Y(_109_));
 OA211x2_ASAP7_75t_SL _236_ (.A1(_118_),
    .A2(_108_),
    .B(_109_),
    .C(net11),
    .Y(_043_));
 INVx1_ASAP7_75t_SL _237_ (.A(\data_in_latch.data_8b_out[6] ),
    .Y(_110_));
 AO21x1_ASAP7_75t_SL _238_ (.A1(_110_),
    .A2(\data_in_latch.data_8b_out[7] ),
    .B(\data_in_latch.data_8b_out[5] ),
    .Y(_111_));
 NAND2x1_ASAP7_75t_SL _239_ (.A(net1),
    .B(_111_),
    .Y(_112_));
 OA211x2_ASAP7_75t_SL _240_ (.A1(net1),
    .A2(_128_),
    .B(_112_),
    .C(net11),
    .Y(_044_));
 NOR2x1_ASAP7_75t_SL _241_ (.A(net1),
    .B(_011_),
    .Y(_113_));
 AND3x1_ASAP7_75t_SL _242_ (.A(\data_in_latch.data_8b_out[5] ),
    .B(_110_),
    .C(net1),
    .Y(_114_));
 OA21x2_ASAP7_75t_SL _243_ (.A1(_113_),
    .A2(_114_),
    .B(net11),
    .Y(_045_));
 INVx1_ASAP7_75t_SL _244_ (.A(_014_),
    .Y(_115_));
 AND3x1_ASAP7_75t_SL _245_ (.A(net11),
    .B(net2),
    .C(_115_),
    .Y(_046_));
 DLLx3_ASAP7_75t_SL _246_ (.CLK(_008_),
    .D(_000_),
    .Q(\data_in_latch.data_8b_out[0] ));
 DLLx3_ASAP7_75t_SL _247_ (.CLK(_008_),
    .D(_001_),
    .Q(\data_in_latch.data_8b_out[1] ));
 DLLx3_ASAP7_75t_SL _248_ (.CLK(_008_),
    .D(_002_),
    .Q(\data_in_latch.data_8b_out[2] ));
 DLLx3_ASAP7_75t_SL _249_ (.CLK(_008_),
    .D(_003_),
    .Q(\data_in_latch.data_8b_out[3] ));
 DLLx3_ASAP7_75t_SL _250_ (.CLK(_008_),
    .D(_004_),
    .Q(\data_in_latch.data_8b_out[4] ));
 DLLx1_ASAP7_75t_SL _251_ (.CLK(_008_),
    .D(_005_),
    .Q(\data_in_latch.data_8b_out[5] ));
 DLLx1_ASAP7_75t_SL _252_ (.CLK(_008_),
    .D(_006_),
    .Q(\data_in_latch.data_8b_out[6] ));
 DLLx1_ASAP7_75t_SL _253_ (.CLK(_008_),
    .D(_007_),
    .Q(\data_in_latch.data_8b_out[7] ));
 DFFLQNx2_ASAP7_75t_SL _254_ (.QN(_027_),
    .CLK(net31),
    .D(_029_));
 DFFLQNx2_ASAP7_75t_SL _255_ (.QN(_026_),
    .CLK(net30),
    .D(_030_));
 DFFLQNx1_ASAP7_75t_SL _256_ (.CLK(net29),
    .D(_031_),
    .QN(_025_));
 DFFLQNx2_ASAP7_75t_SL _257_ (.QN(_024_),
    .CLK(net28),
    .D(_032_));
 DFFLQNx1_ASAP7_75t_SL _258_ (.CLK(net27),
    .D(_033_),
    .QN(_023_));
 DFFLQNx1_ASAP7_75t_SL _259_ (.CLK(net26),
    .D(_034_),
    .QN(_022_));
 DFFLQNx1_ASAP7_75t_SL _260_ (.CLK(net25),
    .D(_035_),
    .QN(_021_));
 DFFLQNx2_ASAP7_75t_SL _261_ (.QN(_020_),
    .CLK(net24),
    .D(_036_));
 DFFLQNx2_ASAP7_75t_SL _262_ (.QN(_019_),
    .CLK(net23),
    .D(_037_));
 DFFLQNx2_ASAP7_75t_SL _263_ (.QN(_018_),
    .CLK(net22),
    .D(_038_));
 DFFLQNx2_ASAP7_75t_SL _264_ (.QN(_017_),
    .CLK(net21),
    .D(_039_));
 DFFLQNx2_ASAP7_75t_SL _265_ (.QN(_016_),
    .CLK(net20),
    .D(_040_));
 DFFLQNx2_ASAP7_75t_SL _266_ (.QN(_015_),
    .CLK(net19),
    .D(_041_));
 DFFLQNx1_ASAP7_75t_SL _267_ (.CLK(net18),
    .D(_042_),
    .QN(_014_));
 DFFLQNx1_ASAP7_75t_SL _268_ (.CLK(net17),
    .D(_043_),
    .QN(_013_));
 DFFLQNx2_ASAP7_75t_SL _269_ (.QN(_012_),
    .CLK(net16),
    .D(_044_));
 DFFLQNx1_ASAP7_75t_SL _270_ (.CLK(net15),
    .D(_045_),
    .QN(_011_));
 DFFLQNx1_ASAP7_75t_SL _271_ (.CLK(net14),
    .D(_046_),
    .QN(_010_));
 DFFLQNx1_ASAP7_75t_SL _272_ (.CLK(net13),
    .D(_047_),
    .QN(_009_));
 TAPCELL_ASAP7_75t_SL PHY_10 ();
 TAPCELL_ASAP7_75t_SL PHY_11 ();
 TAPCELL_ASAP7_75t_SL PHY_12 ();
 TAPCELL_ASAP7_75t_SL PHY_13 ();
 TAPCELL_ASAP7_75t_SL PHY_14 ();
 TAPCELL_ASAP7_75t_SL PHY_15 ();
 TAPCELL_ASAP7_75t_SL PHY_16 ();
 TAPCELL_ASAP7_75t_SL PHY_17 ();
 TAPCELL_ASAP7_75t_SL PHY_18 ();
 TAPCELL_ASAP7_75t_SL PHY_19 ();
 TAPCELL_ASAP7_75t_SL PHY_20 ();
 TAPCELL_ASAP7_75t_SL PHY_21 ();
 TAPCELL_ASAP7_75t_SL PHY_22 ();
 TAPCELL_ASAP7_75t_SL PHY_23 ();
 TAPCELL_ASAP7_75t_SL PHY_24 ();
 TAPCELL_ASAP7_75t_SL PHY_25 ();
 TAPCELL_ASAP7_75t_SL PHY_26 ();
 TAPCELL_ASAP7_75t_SL PHY_27 ();
 TAPCELL_ASAP7_75t_SL PHY_28 ();
 TAPCELL_ASAP7_75t_SL PHY_29 ();
 TAPCELL_ASAP7_75t_SL PHY_30 ();
 TAPCELL_ASAP7_75t_SL PHY_31 ();
 TAPCELL_ASAP7_75t_SL PHY_32 ();
 TAPCELL_ASAP7_75t_SL PHY_33 ();
 TAPCELL_ASAP7_75t_SL PHY_34 ();
 TAPCELL_ASAP7_75t_SL PHY_35 ();
 TAPCELL_ASAP7_75t_SL PHY_36 ();
 TAPCELL_ASAP7_75t_SL PHY_37 ();
 TAPCELL_ASAP7_75t_SL PHY_38 ();
 TAPCELL_ASAP7_75t_SL PHY_39 ();
 TAPCELL_ASAP7_75t_SL PHY_40 ();
 TAPCELL_ASAP7_75t_SL PHY_41 ();
 TAPCELL_ASAP7_75t_SL PHY_42 ();
 TAPCELL_ASAP7_75t_SL PHY_43 ();
 TAPCELL_ASAP7_75t_SL PHY_44 ();
 TAPCELL_ASAP7_75t_SL PHY_45 ();
 TAPCELL_ASAP7_75t_SL PHY_46 ();
 TAPCELL_ASAP7_75t_SL PHY_47 ();
 TAPCELL_ASAP7_75t_SL PHY_48 ();
 TAPCELL_ASAP7_75t_SL PHY_49 ();
 TAPCELL_ASAP7_75t_SL PHY_50 ();
 TAPCELL_ASAP7_75t_SL PHY_51 ();
 TAPCELL_ASAP7_75t_SL PHY_52 ();
 TAPCELL_ASAP7_75t_SL PHY_53 ();
 TAPCELL_ASAP7_75t_SL PHY_54 ();
 TAPCELL_ASAP7_75t_SL PHY_55 ();
 BUFx3_ASAP7_75t_SL input1 (.A(data_en),
    .Y(net1));
 BUFx4f_ASAP7_75t_SL input2 (.A(load_en),
    .Y(net2));
 BUFx2_ASAP7_75t_SL input3 (.A(parallel_data_in[0]),
    .Y(net3));
 BUFx2_ASAP7_75t_SL input4 (.A(parallel_data_in[1]),
    .Y(net4));
 BUFx2_ASAP7_75t_SL input5 (.A(parallel_data_in[2]),
    .Y(net5));
 BUFx2_ASAP7_75t_SL input6 (.A(parallel_data_in[3]),
    .Y(net6));
 BUFx2_ASAP7_75t_SL input7 (.A(parallel_data_in[4]),
    .Y(net7));
 BUFx2_ASAP7_75t_SL input8 (.A(parallel_data_in[5]),
    .Y(net8));
 BUFx2_ASAP7_75t_SL input9 (.A(parallel_data_in[6]),
    .Y(net9));
 BUFx2_ASAP7_75t_SL input10 (.A(parallel_data_in[7]),
    .Y(net10));
 BUFx10_ASAP7_75t_SL input11 (.A(rst_n),
    .Y(net11));
 BUFx2_ASAP7_75t_SL output12 (.A(net12),
    .Y(ser_out));
 INVx1_ASAP7_75t_SL _144__1 (.A(clknet_1_1__leaf_clk),
    .Y(net13));
 INVx1_ASAP7_75t_SL _144__2 (.A(clknet_1_0__leaf_clk),
    .Y(net14));
 INVx1_ASAP7_75t_SL _144__3 (.A(clknet_1_1__leaf_clk),
    .Y(net15));
 INVx1_ASAP7_75t_SL _144__4 (.A(clknet_1_1__leaf_clk),
    .Y(net16));
 INVx1_ASAP7_75t_SL _144__5 (.A(clknet_1_1__leaf_clk),
    .Y(net17));
 INVx1_ASAP7_75t_SL _144__6 (.A(clknet_1_0__leaf_clk),
    .Y(net18));
 INVx1_ASAP7_75t_SL _144__7 (.A(clknet_1_0__leaf_clk),
    .Y(net19));
 INVx1_ASAP7_75t_SL _144__8 (.A(clknet_1_0__leaf_clk),
    .Y(net20));
 INVx1_ASAP7_75t_SL _144__9 (.A(clknet_1_0__leaf_clk),
    .Y(net21));
 INVx1_ASAP7_75t_SL _144__10 (.A(clknet_1_0__leaf_clk),
    .Y(net22));
 INVx1_ASAP7_75t_SL _144__11 (.A(clknet_1_0__leaf_clk),
    .Y(net23));
 INVx1_ASAP7_75t_SL _144__12 (.A(clknet_1_0__leaf_clk),
    .Y(net24));
 INVx1_ASAP7_75t_SL _144__13 (.A(clknet_1_1__leaf_clk),
    .Y(net25));
 INVx1_ASAP7_75t_SL _144__14 (.A(clknet_1_0__leaf_clk),
    .Y(net26));
 INVx1_ASAP7_75t_SL _144__15 (.A(clknet_1_0__leaf_clk),
    .Y(net27));
 INVx1_ASAP7_75t_SL _144__16 (.A(clknet_1_1__leaf_clk),
    .Y(net28));
 INVx1_ASAP7_75t_SL _144__17 (.A(clknet_1_1__leaf_clk),
    .Y(net29));
 INVx1_ASAP7_75t_SL _144__18 (.A(clknet_1_1__leaf_clk),
    .Y(net30));
 INVx1_ASAP7_75t_SL _144__19 (.A(clknet_1_1__leaf_clk),
    .Y(net31));
 BUFx4_ASAP7_75t_SL clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Y(clknet_1_0__leaf_clk));
 BUFx4_ASAP7_75t_SL clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Y(clknet_1_1__leaf_clk));
 DECAPx10_ASAP7_75t_SL FILLER_0_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_0_112 ();
 DECAPx2_ASAP7_75t_SL FILLER_0_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_1_112 ();
 DECAPx2_ASAP7_75t_SL FILLER_1_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_46 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_2_112 ();
 DECAPx2_ASAP7_75t_SL FILLER_2_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_24 ();
 DECAPx1_ASAP7_75t_SL FILLER_3_46 ();
 FILLERxp5_ASAP7_75t_SL FILLER_3_50 ();
 FILLER_ASAP7_75t_SL FILLER_3_55 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_63 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_85 ();
 DECAPx10_ASAP7_75t_SL FILLER_3_107 ();
 DECAPx4_ASAP7_75t_SL FILLER_3_129 ();
 FILLERxp5_ASAP7_75t_SL FILLER_3_139 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_2 ();
 DECAPx6_ASAP7_75t_SL FILLER_4_24 ();
 FILLERxp5_ASAP7_75t_SL FILLER_4_38 ();
 FILLER_ASAP7_75t_SL FILLER_4_42 ();
 FILLER_ASAP7_75t_SL FILLER_4_50 ();
 FILLER_ASAP7_75t_SL FILLER_4_60 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_4_112 ();
 DECAPx2_ASAP7_75t_SL FILLER_4_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_2 ();
 DECAPx6_ASAP7_75t_SL FILLER_5_24 ();
 DECAPx1_ASAP7_75t_SL FILLER_5_38 ();
 FILLERxp5_ASAP7_75t_SL FILLER_5_42 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_5_49 ();
 DECAPx1_ASAP7_75t_SL FILLER_5_59 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_69 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_91 ();
 DECAPx10_ASAP7_75t_SL FILLER_5_113 ();
 DECAPx1_ASAP7_75t_SL FILLER_5_135 ();
 FILLERxp5_ASAP7_75t_SL FILLER_5_139 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_2 ();
 DECAPx2_ASAP7_75t_SL FILLER_6_24 ();
 FILLER_ASAP7_75t_SL FILLER_6_30 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_6_38 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_6_47 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_6_56 ();
 FILLER_ASAP7_75t_SL FILLER_6_71 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_76 ();
 DECAPx10_ASAP7_75t_SL FILLER_6_98 ();
 DECAPx6_ASAP7_75t_SL FILLER_6_120 ();
 DECAPx2_ASAP7_75t_SL FILLER_6_134 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_2 ();
 DECAPx2_ASAP7_75t_SL FILLER_7_24 ();
 FILLERxp5_ASAP7_75t_SL FILLER_7_30 ();
 FILLER_ASAP7_75t_SL FILLER_7_37 ();
 FILLER_ASAP7_75t_SL FILLER_7_46 ();
 DECAPx1_ASAP7_75t_SL FILLER_7_51 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_61 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_83 ();
 DECAPx10_ASAP7_75t_SL FILLER_7_105 ();
 DECAPx4_ASAP7_75t_SL FILLER_7_127 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_7_137 ();
 DECAPx1_ASAP7_75t_SL FILLER_8_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_11 ();
 DECAPx2_ASAP7_75t_SL FILLER_8_33 ();
 FILLERxp5_ASAP7_75t_SL FILLER_8_39 ();
 DECAPx1_ASAP7_75t_SL FILLER_8_46 ();
 FILLERxp5_ASAP7_75t_SL FILLER_8_50 ();
 DECAPx1_ASAP7_75t_SL FILLER_8_57 ();
 FILLERxp5_ASAP7_75t_SL FILLER_8_61 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_68 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_90 ();
 DECAPx10_ASAP7_75t_SL FILLER_8_112 ();
 DECAPx2_ASAP7_75t_SL FILLER_8_134 ();
 DECAPx4_ASAP7_75t_SL FILLER_9_2 ();
 FILLER_ASAP7_75t_SL FILLER_9_12 ();
 DECAPx4_ASAP7_75t_SL FILLER_9_20 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_9_30 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_9_39 ();
 FILLER_ASAP7_75t_SL FILLER_9_49 ();
 FILLER_ASAP7_75t_SL FILLER_9_57 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_69 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_9_91 ();
 FILLER_ASAP7_75t_SL FILLER_9_102 ();
 DECAPx10_ASAP7_75t_SL FILLER_9_110 ();
 DECAPx2_ASAP7_75t_SL FILLER_9_132 ();
 FILLER_ASAP7_75t_SL FILLER_9_138 ();
 DECAPx1_ASAP7_75t_SL FILLER_10_2 ();
 FILLER_ASAP7_75t_SL FILLER_10_11 ();
 DECAPx1_ASAP7_75t_SL FILLER_10_30 ();
 FILLER_ASAP7_75t_SL FILLER_10_39 ();
 DECAPx2_ASAP7_75t_SL FILLER_10_50 ();
 DECAPx4_ASAP7_75t_SL FILLER_10_62 ();
 DECAPx4_ASAP7_75t_SL FILLER_10_80 ();
 DECAPx2_ASAP7_75t_SL FILLER_10_93 ();
 FILLERxp5_ASAP7_75t_SL FILLER_10_99 ();
 FILLER_ASAP7_75t_SL FILLER_10_108 ();
 DECAPx10_ASAP7_75t_SL FILLER_10_116 ();
 FILLER_ASAP7_75t_SL FILLER_10_138 ();
 DECAPx2_ASAP7_75t_SL FILLER_11_2 ();
 FILLER_ASAP7_75t_SL FILLER_11_8 ();
 FILLER_ASAP7_75t_SL FILLER_11_16 ();
 DECAPx2_ASAP7_75t_SL FILLER_11_35 ();
 FILLER_ASAP7_75t_SL FILLER_11_41 ();
 FILLER_ASAP7_75t_SL FILLER_11_49 ();
 DECAPx1_ASAP7_75t_SL FILLER_11_61 ();
 DECAPx6_ASAP7_75t_SL FILLER_11_73 ();
 FILLER_ASAP7_75t_SL FILLER_11_87 ();
 FILLER_ASAP7_75t_SL FILLER_11_97 ();
 DECAPx1_ASAP7_75t_SL FILLER_11_102 ();
 FILLERxp5_ASAP7_75t_SL FILLER_11_106 ();
 DECAPx10_ASAP7_75t_SL FILLER_11_113 ();
 DECAPx1_ASAP7_75t_SL FILLER_11_135 ();
 FILLERxp5_ASAP7_75t_SL FILLER_11_139 ();
 DECAPx1_ASAP7_75t_SL FILLER_12_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_11 ();
 DECAPx2_ASAP7_75t_SL FILLER_12_33 ();
 FILLERxp5_ASAP7_75t_SL FILLER_12_39 ();
 DECAPx2_ASAP7_75t_SL FILLER_12_46 ();
 FILLER_ASAP7_75t_SL FILLER_12_55 ();
 DECAPx2_ASAP7_75t_SL FILLER_12_64 ();
 FILLER_ASAP7_75t_SL FILLER_12_70 ();
 DECAPx2_ASAP7_75t_SL FILLER_12_81 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_12_87 ();
 DECAPx2_ASAP7_75t_SL FILLER_12_93 ();
 FILLER_ASAP7_75t_SL FILLER_12_99 ();
 FILLER_ASAP7_75t_SL FILLER_12_109 ();
 DECAPx10_ASAP7_75t_SL FILLER_12_117 ();
 FILLERxp5_ASAP7_75t_SL FILLER_12_139 ();
 FILLER_ASAP7_75t_SL FILLER_13_2 ();
 FILLER_ASAP7_75t_SL FILLER_13_9 ();
 FILLER_ASAP7_75t_SL FILLER_13_17 ();
 FILLER_ASAP7_75t_SL FILLER_13_36 ();
 DECAPx2_ASAP7_75t_SL FILLER_13_44 ();
 FILLER_ASAP7_75t_SL FILLER_13_50 ();
 DECAPx1_ASAP7_75t_SL FILLER_13_59 ();
 FILLER_ASAP7_75t_SL FILLER_13_69 ();
 DECAPx4_ASAP7_75t_SL FILLER_13_79 ();
 FILLER_ASAP7_75t_SL FILLER_13_92 ();
 FILLER_ASAP7_75t_SL FILLER_13_97 ();
 DECAPx2_ASAP7_75t_SL FILLER_13_107 ();
 DECAPx6_ASAP7_75t_SL FILLER_13_119 ();
 DECAPx2_ASAP7_75t_SL FILLER_13_133 ();
 FILLERxp5_ASAP7_75t_SL FILLER_13_139 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_2 ();
 DECAPx4_ASAP7_75t_SL FILLER_14_24 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_14_34 ();
 FILLER_ASAP7_75t_SL FILLER_14_43 ();
 FILLER_ASAP7_75t_SL FILLER_14_51 ();
 DECAPx6_ASAP7_75t_SL FILLER_14_60 ();
 FILLERxp5_ASAP7_75t_SL FILLER_14_74 ();
 DECAPx4_ASAP7_75t_SL FILLER_14_78 ();
 FILLER_ASAP7_75t_SL FILLER_14_88 ();
 DECAPx10_ASAP7_75t_SL FILLER_14_110 ();
 DECAPx2_ASAP7_75t_SL FILLER_14_132 ();
 FILLER_ASAP7_75t_SL FILLER_14_138 ();
 DECAPx2_ASAP7_75t_SL FILLER_15_2 ();
 DECAPx1_ASAP7_75t_SL FILLER_15_14 ();
 FILLERxp5_ASAP7_75t_SL FILLER_15_18 ();
 FILLER_ASAP7_75t_SL FILLER_15_36 ();
 DECAPx1_ASAP7_75t_SL FILLER_15_47 ();
 FILLERxp5_ASAP7_75t_SL FILLER_15_51 ();
 DECAPx4_ASAP7_75t_SL FILLER_15_60 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_15_70 ();
 DECAPx1_ASAP7_75t_SL FILLER_15_94 ();
 FILLERxp5_ASAP7_75t_SL FILLER_15_98 ();
 FILLER_ASAP7_75t_SL FILLER_15_120 ();
 DECAPx6_ASAP7_75t_SL FILLER_15_125 ();
 FILLERxp5_ASAP7_75t_SL FILLER_15_139 ();
 DECAPx6_ASAP7_75t_SL FILLER_16_2 ();
 FILLERxp5_ASAP7_75t_SL FILLER_16_16 ();
 DECAPx4_ASAP7_75t_SL FILLER_16_34 ();
 DECAPx2_ASAP7_75t_SL FILLER_16_50 ();
 FILLERxp5_ASAP7_75t_SL FILLER_16_56 ();
 FILLER_ASAP7_75t_SL FILLER_16_65 ();
 FILLER_ASAP7_75t_SL FILLER_16_73 ();
 FILLER_ASAP7_75t_SL FILLER_16_96 ();
 FILLER_ASAP7_75t_SL FILLER_16_101 ();
 DECAPx1_ASAP7_75t_SL FILLER_16_106 ();
 FILLER_ASAP7_75t_SL FILLER_16_116 ();
 DECAPx6_ASAP7_75t_SL FILLER_16_124 ();
 FILLER_ASAP7_75t_SL FILLER_16_138 ();
 FILLER_ASAP7_75t_SL FILLER_17_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_17_9 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_18 ();
 DECAPx10_ASAP7_75t_SL FILLER_17_40 ();
 DECAPx2_ASAP7_75t_SL FILLER_17_62 ();
 FILLER_ASAP7_75t_SL FILLER_17_68 ();
 FILLER_ASAP7_75t_SL FILLER_17_73 ();
 FILLER_ASAP7_75t_SL FILLER_17_96 ();
 FILLER_ASAP7_75t_SL FILLER_17_118 ();
 FILLER_ASAP7_75t_SL FILLER_17_128 ();
 FILLER_ASAP7_75t_SL FILLER_17_138 ();
 DECAPx2_ASAP7_75t_SL FILLER_18_2 ();
 FILLER_ASAP7_75t_SL FILLER_18_8 ();
 DECAPx10_ASAP7_75t_SL FILLER_18_16 ();
 DECAPx6_ASAP7_75t_SL FILLER_18_38 ();
 DECAPx1_ASAP7_75t_SL FILLER_18_52 ();
 FILLERxp5_ASAP7_75t_SL FILLER_18_56 ();
 FILLER_ASAP7_75t_SL FILLER_18_67 ();
 FILLER_ASAP7_75t_SL FILLER_18_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_18_99 ();
 DECAPx6_ASAP7_75t_SL FILLER_18_122 ();
 DECAPx1_ASAP7_75t_SL FILLER_18_136 ();
 FILLER_ASAP7_75t_SL FILLER_19_2 ();
 FILLER_ASAP7_75t_SL FILLER_19_9 ();
 DECAPx1_ASAP7_75t_SL FILLER_19_16 ();
 FILLERxp5_ASAP7_75t_SL FILLER_19_20 ();
 FILLER_ASAP7_75t_SL FILLER_19_27 ();
 DECAPx4_ASAP7_75t_SL FILLER_19_44 ();
 DECAPx2_ASAP7_75t_SL FILLER_19_58 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_19_64 ();
 FILLER_ASAP7_75t_SL FILLER_19_70 ();
 FILLER_ASAP7_75t_SL FILLER_19_75 ();
 FILLER_ASAP7_75t_SL FILLER_19_98 ();
 FILLER_ASAP7_75t_SL FILLER_19_103 ();
 DECAPx2_ASAP7_75t_SL FILLER_19_125 ();
 FILLER_ASAP7_75t_SL FILLER_19_131 ();
 FILLER_ASAP7_75t_SL FILLER_19_138 ();
 DECAPx2_ASAP7_75t_SL FILLER_20_2 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_20_8 ();
 DECAPx4_ASAP7_75t_SL FILLER_20_26 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_20_36 ();
 DECAPx10_ASAP7_75t_SL FILLER_20_42 ();
 DECAPx6_ASAP7_75t_SL FILLER_20_64 ();
 FILLERxp5_ASAP7_75t_SL FILLER_20_78 ();
 DECAPx4_ASAP7_75t_SL FILLER_20_82 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_20_92 ();
 FILLER_ASAP7_75t_SL FILLER_20_115 ();
 FILLER_ASAP7_75t_SL FILLER_20_120 ();
 FILLER_ASAP7_75t_SL FILLER_20_125 ();
 DECAPx4_ASAP7_75t_SL FILLER_20_130 ();
 FILLER_ASAP7_75t_SL FILLER_21_2 ();
 FILLER_ASAP7_75t_SL FILLER_21_9 ();
 DECAPx2_ASAP7_75t_SL FILLER_21_26 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_21_32 ();
 FILLER_ASAP7_75t_SL FILLER_21_47 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_21_55 ();
 DECAPx2_ASAP7_75t_SL FILLER_21_78 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_21_84 ();
 FILLER_ASAP7_75t_SL FILLER_21_90 ();
 FILLER_ASAP7_75t_SL FILLER_21_99 ();
 DECAPx2_ASAP7_75t_SL FILLER_21_121 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_21_127 ();
 DECAPx2_ASAP7_75t_SL FILLER_21_133 ();
 FILLERxp5_ASAP7_75t_SL FILLER_21_139 ();
 DECAPx2_ASAP7_75t_SL FILLER_22_2 ();
 FILLER_ASAP7_75t_SL FILLER_22_8 ();
 DECAPx6_ASAP7_75t_SL FILLER_22_16 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_22_30 ();
 FILLER_ASAP7_75t_SL FILLER_22_39 ();
 FILLER_ASAP7_75t_SL FILLER_22_47 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_22_57 ();
 DECAPx2_ASAP7_75t_SL FILLER_22_67 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_22_73 ();
 DECAPx4_ASAP7_75t_SL FILLER_22_79 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_22_89 ();
 DECAPx1_ASAP7_75t_SL FILLER_22_99 ();
 FILLERxp5_ASAP7_75t_SL FILLER_22_103 ();
 FILLER_ASAP7_75t_SL FILLER_22_110 ();
 FILLER_ASAP7_75t_SL FILLER_22_120 ();
 DECAPx6_ASAP7_75t_SL FILLER_22_125 ();
 FILLERxp5_ASAP7_75t_SL FILLER_22_139 ();
 FILLER_ASAP7_75t_SL FILLER_23_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_23_18 ();
 DECAPx2_ASAP7_75t_SL FILLER_23_40 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_23_46 ();
 DECAPx1_ASAP7_75t_SL FILLER_23_55 ();
 FILLERxp5_ASAP7_75t_SL FILLER_23_59 ();
 DECAPx1_ASAP7_75t_SL FILLER_23_66 ();
 FILLERxp5_ASAP7_75t_SL FILLER_23_70 ();
 FILLER_ASAP7_75t_SL FILLER_23_91 ();
 FILLER_ASAP7_75t_SL FILLER_23_115 ();
 FILLER_ASAP7_75t_SL FILLER_23_138 ();
 DECAPx10_ASAP7_75t_SL FILLER_24_2 ();
 DECAPx6_ASAP7_75t_SL FILLER_24_24 ();
 DECAPx2_ASAP7_75t_SL FILLER_24_38 ();
 FILLERxp5_ASAP7_75t_SL FILLER_24_44 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_24_51 ();
 FILLER_ASAP7_75t_SL FILLER_24_60 ();
 FILLER_ASAP7_75t_SL FILLER_24_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_24_91 ();
 FILLER_ASAP7_75t_SL FILLER_24_115 ();
 FILLER_ASAP7_75t_SL FILLER_24_120 ();
 DECAPx4_ASAP7_75t_SL FILLER_24_129 ();
 FILLERxp5_ASAP7_75t_SL FILLER_24_139 ();
 DECAPx10_ASAP7_75t_SL FILLER_25_2 ();
 DECAPx6_ASAP7_75t_SL FILLER_25_24 ();
 DECAPx1_ASAP7_75t_SL FILLER_25_38 ();
 FILLERxp5_ASAP7_75t_SL FILLER_25_42 ();
 DECAPx2_ASAP7_75t_SL FILLER_25_51 ();
 FILLERxp5_ASAP7_75t_SL FILLER_25_57 ();
 FILLER_ASAP7_75t_SL FILLER_25_66 ();
 DECAPx1_ASAP7_75t_SL FILLER_25_76 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_SL FILLER_25_100 ();
 DECAPx1_ASAP7_75t_SL FILLER_25_109 ();
 FILLER_ASAP7_75t_SL FILLER_25_119 ();
 FILLER_ASAP7_75t_SL FILLER_25_124 ();
 DECAPx4_ASAP7_75t_SL FILLER_25_129 ();
 FILLERxp5_ASAP7_75t_SL FILLER_25_139 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_24 ();
 DECAPx6_ASAP7_75t_SL FILLER_26_46 ();
 FILLER_ASAP7_75t_SL FILLER_26_60 ();
 FILLER_ASAP7_75t_SL FILLER_26_65 ();
 FILLER_ASAP7_75t_SL FILLER_26_70 ();
 FILLER_ASAP7_75t_SL FILLER_26_93 ();
 FILLER_ASAP7_75t_SL FILLER_26_98 ();
 DECAPx10_ASAP7_75t_SL FILLER_26_103 ();
 DECAPx6_ASAP7_75t_SL FILLER_26_125 ();
 FILLERxp5_ASAP7_75t_SL FILLER_26_139 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_2 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_24 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_46 ();
 DECAPx2_ASAP7_75t_SL FILLER_27_68 ();
 FILLER_ASAP7_75t_SL FILLER_27_74 ();
 FILLER_ASAP7_75t_SL FILLER_27_79 ();
 DECAPx1_ASAP7_75t_SL FILLER_27_87 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_94 ();
 DECAPx10_ASAP7_75t_SL FILLER_27_116 ();
 FILLER_ASAP7_75t_SL FILLER_27_138 ();
endmodule
